-- ROM_mem.vhd
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ROM_mem is
    Port (enable : in std_logic;
          h_pos : in std_logic_vector(9 downto 0);
          v_pos : in std_logic_vector(9 downto 0);
          data : out std_logic_vector(3 downto 0));
end ROM_mem;

architecture Behavioral of ROM_mem is
type rom_type is array(0 to 479, 0 to 639) of std_logic_vector(3 downto 0); -- 640x480 image resolution
--type rom_type is array(0 to 66, 0 to 99) of std_logic_vector(3 downto 0); -- 100x67 image resolution
   -- ROM image:
constant ROM: rom_type :=(
("0111","0111","0111","0111","0111","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1011","1010","1010","1010","1010","1011","1010","1010","1011","1011","1011","1011","1011","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1011","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001"),
("0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","1011","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001"),
("1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1000","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1010","1010","1010","1010","1011","1011","1011","1010","1011","1011","1011","1011","1010","1010","1010","1011","1011","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1010","1011","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","1011","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1000","1001","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1000","1001","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1010","1010","1011","1011","1011","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1011","1011","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1010","1001","1010","1001","1010","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1010","1010","1010","1010","1010","1001","1010","1001","1010","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1000","1000","1001","1001","1000","1000"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1001","1001","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1001","1000","1001"),
("1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1001","1010","1001","1001","1001","1010","1010","1010","1001","1001","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1001","1001","1001","1000","1000","1001","1001","1000","1000","1001","1000","1001","1001","1001"),
("1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000"),
("1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1010","1010","1010","1001","1001","1001","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1000","1001","1000","1000","1000","1001","1001","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1001","1001","1010","1010","1001","1010","1010","1001","1010","1001","1001","1001","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1001","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1010","1010","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1001","1000","1001","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1010","1001","1010","1010","1010","1001","1010","1001","1010","1001","1001","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1001","1010","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1001","1001","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1010","1010","1010","1010","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1010","1010","1010","1010","1010","1011","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1001","1001","1001","1001","1001","1000","1001","1000","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","1000","0111","1000","0111","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1010","1010","1010","1011","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1011","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1000","1000","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","1000","0111","1000","0111","1000","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1001","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1011","1010","1011","1011","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1001","1001","1000","1000","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1001","1001","1001","1010","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1001","1010","1010","1010","1001","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1010","1010","1010","1011","1011","1011","1011","1010","1011","1011","1011","1010","1011","1011","1011","1011","1011","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1010","1011","1011","1010","1011","1011","1011","1011","1011","1010","1010","1011","1011","1010","1010","1010","1011","1011","1011","1010","1010","1010","1011","1011","1010","1011","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1001","1010","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1001","1001","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1011","1010","1010","1010","1011","1011","1011","1010","1010","1010","1010","1011","1010","1011","1010","1010","1011","1011","1011","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1010","1010","1001","1010","1010","1001","1001","1001","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1011","1010","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1010","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","0111","1000","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1010","1001","1010","1001","1001","1010","1010","1001","1001","1010","1010","1010","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1011","1011","1010","1010","1011","1010","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1010","1010","1001","1010","1001","1010","1001","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1001","1010","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1001","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1011","1010","1011","1011","1010","1010","1010","1011","1010","1011","1011","1011","1011","1011","1011","1010","1011","1010","1011","1011","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1011","1010","1011","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1001","1001","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1010","1010","1010","1011","1010","1010","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1001","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1011","1011","1010","1011","1011","1011","1010","1011","1011","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1011","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","0111","0111","1000","1000","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1011","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1011","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1010","1011","1010","1010","1010","1011","1011","1011","1010","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","0111","1000","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1010","1010","1010","1011","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","1011","1011","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1000","1001","1000","1000","1001","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1011","1010","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1010","1011","1011","1010","1011","1010","1010","1011","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1010","1010","1010","1010","1010","1011","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1010","1010","1011","1010","1010","1010","1011","1011","1011","1010","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1001","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","1000","0111","1000","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1011","1011","1010","1010","1011","1011","1010","1010","1010","1011","1011","1010","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1010","1010","1011","1011","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1001","1001","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","1011","1011","1010","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1001","1001","1000","1000","1001","1001","1001","1001","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1010","1011","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1010","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1000","1000","1000","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1010","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1011","1010","1010","1011","1011","1010","1011","1010","1010","1010","1011","1011","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1001","1000","1001","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0111","0111","0111","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","1000","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1011","1010","1011","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1000","1000","1000","1001","1000","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0111","0110","0110","0110","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1011","1010","1010","1011","1010","1011","1011","1010","1011","1010","1011","1011","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1001","1001","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1011","1010","1010","1010","1010","1011","1010","1011","1011","1011","1011","1011","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1011","1010","1011","1010","1010","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1010","1010","1010","1011","1011","1011","1011","1011","1010","1011","1011","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1001","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1010","1010","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","1010","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1001","1010","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0111","0110","0111","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1010","1010","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1001","1001","1001","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","1010","1011","1011","1010","1011","1010","1010","1011","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1010","1010","1010","1011","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1010","1001","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1001","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1010","1011","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1001","1010","1010","1001","1001","1010","1001","1001","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1001","1010","1001","1001","1010","1001","1010","1010","1010","1001","1001","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1001","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1011","1011","1011","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1010","1010","1011","1011","1011","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000"),
("0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0111","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1001","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1010","1011","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","0111"),
("0110","0110","0111","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1010","1011","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000"),
("0110","0110","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1010","1011","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1010","1010","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1011","1011","1011","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1011","1011","1010","1010","1010","1011","1011","1011","1011","1010","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1010","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","1011","1010","1010","1011","1010","1010","1011","1011","1010","1011","1011","1011","1011","1010","1011","1011","1011","1011","1010","1011","1011","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1011","1011","1011","1011","1010","1011","1011","1011","1010","1011","1011","1011","1010","1010","1011","1011","1010","1010","1011","1010","1010","1011","1010","1010","1011","1011","1011","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1011","1011","1011","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1001","1001","1010","1001","1010","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1000","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1011","1010","1011","1011","1011","1010","1011","1010","1010","1010","1010","1011","1010","1010","1011","1011","1010","1010","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1011","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1010","1001","1010","1010","1001","1010","1001","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1011","1010","1011","1010","1010","1011","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1000","1000","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1001","1010","1001","1010","1010","1010","1010","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","1000","0111","1000","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1001","1000","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1001","1001","1001","1010","1010","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","1000","0111","1000","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1001","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","0111","0111","0111","0111","1000","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1000","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","1000","0111","1000","0111","1000","1000","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1001","1001","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","0011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1010","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","0111","0111","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","1000","0111","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","0011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1010","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1001","1001","1001","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1001","1001","1001","1010","1010","1010","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0100","0011","0011","0010","0011","0100","0110","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1000","0110","0011","0110","0111","1000","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1001","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0010","1001","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","0100","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","0100","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0100","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","1000","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0100","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1001","1010","1010","1001","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1001","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0100","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1001","1010","1010","1010","1010","1001","1001","1010","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0010","0101","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1000","1000","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0010","0001","0001","0111","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1000","1000","1000","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0100","0000","0000","0000","0100","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1001","1010","1010","1010","1001","1001","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","0110","0000","0101","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0000","0111","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0001","0110","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0111","0000","0110","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0110","0000","0101","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","1000","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0101","0000","0011","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0100","0000","0010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0011","0000","0010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","0010","0001","0001","1000","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1001","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0001","0001","0000","0111","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1000","1001","1000","1000","1001","1001","1001","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0001","0001","0000","0110","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1000","1001","1001","1001","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0110","0001","0001","0001","0101","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1001","1010","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1000","1001","1001","1000","1000","1001","1000","1000","1000","1001","1001","1000","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1010","1001","1001","1001","1001","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0101","0001","0001","0001","0011","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1001","1001","1001","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1010","1010","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0100","0001","0001","0001","0011","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1010","1001","1001","1010","1010","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0011","0001","0010","0001","0010","1000","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","0010","0001","0010","0001","0001","0111","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1010","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0010","0001","0010","0001","0001","0110","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1001","1010","1010","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0001","0010","0010","0010","0001","0101","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1010","1001","1010","1010","1010","1001","1001","1010","1010","1001","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0111","0001","0010","0010","0010","0001","0101","1010","1010","1001","1001","1001","1010","1001","1001","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1010","1010","1001","1001","1010","1001","1010","1010","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1010","1001","1001","1010","1010","1010","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0110","0001","0010","0010","0010","0001","0011","1001","1001","1001","1010","1001","1001","1001","1001","1010","1010","1010","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1001","1010","1010","1010","1001","1010","1001","1010","1010","1001","1001","1001","1010","1001","1010","1010","1001","1010","1010","1010","1001","1010","1010","1010","1001","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","0101","0001","0010","0010","0010","0001","0010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1001","1001","1010","1001","1001","1001","1001","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1010","1001","1010","1010","1010","0100","0001","0010","0010","0010","0001","0010","1000","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1001","1001","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1010","1010","1001","1001","1010","1010","1001","1001","1010","1001","1010","1010","1001","0011","0010","0010","0010","0010","0001","0001","1000","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1010","1010","1001","1001","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1010","1001","1010","1001","0010","0010","0010","0010","0010","0010","0001","0110","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1001","1001","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1001","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1001","1001","1001","1010","1001","1010","1001","1001","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1000","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1010","1001","1001","1001","1001","1010","1010","1001","1001","1010","1001","1010","1010","1010","1010","1001","1010","1001","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1010","1010","1010","1000","0010","0010","0010","0010","0010","0010","0001","0101","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1001","1001","1001","1001","1010","1001","1001","1010","1001","1001","1001","1010","1010","1010","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1000","1001","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1001","1001","1000","1000","1001","1000","1001","1001","1001","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1001","1001","1001","1001","1010","1001","1010","1010","1001","1001","1010","1010","1010","1010","1001","1001","1001","1001","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1010","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1010","1010","1001","1001","1010","1010","1001","1001","1001","1001","1010","1010","0111","0001","0010","0010","0010","0010","0010","0001","0100","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1001","1000","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","1000","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1001","1001","1001","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0110","0001","0010","0010","0010","0010","0010","0001","0011","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1001","1001","1001","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1001","1001","1010","1001","1001","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","0101","0001","0010","0010","0010","0010","0010","0001","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","0111","1000","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1001","1001","1000","1001","1001","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","0100","0001","0010","0010","0010","0010","0010","0010","0010","1000","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1001","1010","1001","1010","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1001","1000","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1010","1010","1010","1001","1010","1001","1001","1001","1001","1010","1010","1001","1001","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","0011","0010","0010","0010","0010","0010","0010","0010","0001","0111","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1001","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1001","1010","1001","1001","1010","1010","1010","1001","1001","1010","1010","1010","1001","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0110","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1001","1001","1001","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1001","1001","1010","1001","1010","1010","1010","1001","1001","1001","1001","1001","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1000","0010","0010","0010","0010","0010","0010","0010","0010","0001","0101","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1001","1001","1010","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1010","1010","1001","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0111","0010","0010","0010","0010","0010","0010","0010","0010","0001","0100","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0110","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1001","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1010","1001","1010","1010","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1000","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1000","1000","1001","1000","1000","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1001","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1010","1001","1010","1001","1010","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0110","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","1000","0111","1000","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1001","1001","1000","1000","1000","1000","1000","1001","1001","1001","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0001","0101","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1000","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0001","0100","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0111","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0001","0011","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","1000","0111","0111","0111","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0110","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0001","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0101","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0100","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1001","1001","1001","1001","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0011","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0110","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0101","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0100","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0111","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1000","1001","1000","1000","1001","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0110","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0101","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0100","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0110","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1001","1001","1001","1001","1000","1000","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0101","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0100","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1000","1001","1000","1000","1000","1001","1000","1000","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1001","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0111","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0110","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0101","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0100","0001","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0100","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","1000","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1001","1001","1000","1000","1001","1001","1000","1001","1001","1001","1001","1000","1000","1001","1001","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1000","0011","0011","0011","0100","0100","0011","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0111"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1000","1001","1000","1000","1001","1000","1001","1000","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","0101","0011","0011","0100","0100","0100","0011","0100","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0010","0100","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0110","0011","0011","0011","0100","0100","0011","0011","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0110","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1000","1001","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1000","0011","0011","0011","0011","0100","0100","0011","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","0111","0111","0111","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1001","1000","1000","1001","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0100","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0110","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0110","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0010","0010","0010","0010","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0110","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0001","0010","0010","0010","0001","0010","0010","0010","0010","0001","0001","0010","0010","0011","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1000","0100","0011","0011","0010","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0001","0011","0011","0100","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1000","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","0101","0101","0101","0011","0100","0101","0101","0110","0100","0100","0100","0100","0101","0101","0101","0110","0110","0110","0101","0100","0011","0100","0100","0101","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1000","1001","1000","1000","1001","1000","1000","1000","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0110","0110","0101","0101","0101","0110","0110","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1000","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1000","1000","1001","1001","1001","1001","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0011","0111","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0100","0110","0100","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1001","1000","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0100","1000","0101","0011","0011","0011","0011","0100","0100","0011","0011","0011","0010","0100","0100","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0100","0111","0100","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1001","1000","1001","1001","1001","1001","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0111","0110","0111","0111","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0100","0111","0101","0011","0011","0011","0011","0100","0100","0100","0100","0011","0010","0100","0100","0011","0011","0100","0100","0011","0011","0100","0100","0100","0011","0100","0110","0100","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1000","1001","1000","1000","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1000","0011","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0100","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1001","1000","1000","1001","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1001","1001","1001","1000","1000","1001","1001","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1000","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0101","0101","0011","0011","0011","0011","0011","0100","0100","0011","0100","0011","0100","0100","0010","1000","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0111","0011","0100","0101","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0101","0101","0011","0011","0011","0100","0100","0100","0011","0100","0100","0011","0101","0100","0010","0111","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110"),
("0111","0110","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0111","0010","0100","0111","0101","0100","0101","0101","0101","0101","0100","0100","0100","0011","0101","0101","0011","0011","0100","0100","0101","0101","0101","0100","0101","0101","0110","0100","0011","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101"),
("0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0111","0011","0011","0101","0101","0110","0110","0110","0110","0110","0101","0100","0100","0100","0110","0110","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0011","0011","0110","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1001","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","1000","1000","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0100"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0100","0010","0001","0011","0101","0110","0110","0110","0110","0101","0101","0100","0100","0010","0010","0010","0010","0011","0100","0101","0110","0101","0101","0110","0101","0101","0100","0001","0001","0011","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","0111","0111","1000","0111","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0100","0100","0101","0101","0101","0100"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0101","0010","0001","0100","0101","0101","0100","0100","0110","0110","0101","0100","0100","0011","0100","0100","0011","0100","0100","0101","0110","0110","0100","0011","0100","0101","0100","0010","0010","0100","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","0111","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0110","0111","0110","0101","0111","0111","0111","0111","0111","0110","0101","0100","0100","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0101","0100","0101","0110","0110","0101","0101","0101","0101","0110","0101","0101","0101","0100","0101","0101","0110","0110","0110","0110","0101","0101","0101"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0011","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0110","0011","0010","0100","0101","0011","0010","0011","0100","0101","0101","0100","0100","0011","0100","0100","0011","0100","0100","0101","0110","0100","0010","0010","0011","0100","0101","0010","0011","0101","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0110","0110","0110","1000","1000","0111","1000","1000","1000","1001","1000","1001","1001","1001","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0101","0110","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0101","0101","0111","0111","0110","0101","0110","0110","0111","1000","0110","0110","0101","0100","0100","0101","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0110","0110","0110","0110","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0100","0100","0100","0100","0100","0100","0110","0111","0101","0110","0111","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0110"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0011","0011","0100","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","0111","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0110","0011","0011","0100","0011","0101","0011","0010","0100","0100","0101","0101","0100","0011","0100","0100","0011","0011","0100","0101","0101","0011","0010","0001","0011","0011","0100","0010","0010","0100","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","0111","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","0111","0110","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0110","0110","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","0110","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0100","0100","0100","0100","0101","0100","0101","0101","0101","0101","0110","0110","0100","0101","0101","0101","0101","0101","0101","0101","0101","0110","0111"),
("0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0010","0011","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0111","0110","0111","0110","0111","0110","0111","0110","0110","0110","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0101","0011","0010","0011","0100","0110","0100","0011","0101","0101","0101","0101","0100","0011","0100","0100","0011","0100","0101","0101","0101","0100","0101","0010","0100","0011","0100","0010","0010","0100","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","0111","1000","1000","1000","0111","0111","0111","0111","1000","1000","0111","1000","1000","1000","0111","1000","1000","1000","0111","0111","0111","0111","1000","1000","1001","1000","1000","1000","1000","0111","1000","0111","1000","1000","0111","1000","0111","0110","0111","1000","0111","0111","1000","0111","1000","1000","1000","1000","1001","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","1000","1000","0111","1000","1000","1000","0111","0111","0111","1000","0111","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","1000","1000","0111","0111","1000","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0110","0111","0110","0110","0110","0111","0110","0111","1000","0111","0110","0111","1000","0110","0110","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0110","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0110","0101","0101","0111","0110","0110","0110","0100","0100","0111"),
("0110","0110","0110","0110","0110","0100","0101","0101","0101","0101","0011","0010","0011","0100","0011","0011","0101","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","1000","1001","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1000","1000","1000","1000","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","1000","1000","1000","0111","0111","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0101","0011","0011","0100","0100","0101","0110","0101","0110","0011","0101","0101","0100","0011","0100","0100","0011","0100","0100","0101","0100","0100","0110","0100","0101","0010","0100","0010","0010","0100","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","0111","0111","0111","1000","0111","1000","0111","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","0111","1000","0111","1000","1001","1001","1001","0110","0100","0101","1001","1001","1001","1001","1000","0111","0111","0111","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0110","0101","0101","0101","0101","0110","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","1000","1000","0110","0110","1000","1000","0110","0111","0110","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0110","0111","0111","1000","1000","0111","0111","0111","1000","0111","0110","0111","0101","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0101","0101","0101","0110","0101","0101","0100","0101","0101","0100","0100","0100","0100","0100","0101","0101","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0110","0110","0101","0111","0111","0111","0111","0111","0110","0111"),
("0110","0110","0110","0111","0110","0010","0110","0111","0111","0101","0010","0001","0001","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","0110","0011","0011","0100","0100","0011","0100","0101","0101","0011","0101","0101","0100","0011","0100","0100","0011","0011","0100","0100","0100","0010","0100","0011","0011","0011","0100","0010","0010","0100","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0101","0101","0110","1000","0111","1000","0111","1000","1000","0111","0111","1001","1001","1001","0110","0100","0101","1001","1001","1001","1001","0111","0110","0110","0111","1000","1000","1000","1000","1000","1000","1001","1000","1000","1001","1001","1000","1000","1000","0111","0111","0111","0111","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","0111","1000","1000","1000","0111","1000","1000","0111","0111","1000","1000","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0110","0110","0110","0111","1000","0111","0111","1000","0111","0111","1000","1000","0111","0111","1000","1000","0111","0111","0111","0111","0110","0101","0101","0101","0101","0101","0110","0110","0101","0110","0111","0110","0111","1000","0111","0110","0111","1000","0110","0110","0111","0101","0100","0101","0101","0100","0101","0101","0110","0110","0110","0110","0101","0110","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0110","0110","0100","0100","0100","0100","0101","0100","0100","0100","0011","0100","0101","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0110","0110","0110","0101","0100","0010","0011","0100","0100","0010","0001","0001","0001","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0111","0110","0111","0110","0110","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","0110","0100","0011","0100","0101","0011","0010","0100","0101","0100","0101","0101","0101","0100","0100","0100","0011","0011","0100","0100","0100","0011","0010","0010","0011","0100","0101","0011","0011","0100","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","1000","1000","1000","1000","0111","0110","0110","0110","0111","0111","0110","1000","1001","1001","1000","0101","0101","0110","1000","1001","1000","0111","1000","1000","0111","0110","1001","1010","1001","0110","0100","0101","1001","1001","1001","1001","0111","0110","0110","0110","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","1000","0111","0111","0111","1000","0111","1000","0111","0111","1000","0111","0111","1000","0111","1000","1000","1000","0111","1000","0111","0111","0111","0111","1000","0111","0111","0111","1000","0111","1000","0111","0111","1000","1000","1000","1000","0111","1000","1000","1000","0111","1000","0111","0111","0110","0101","0101","0110","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0101","0101","0101","0110","0110","0110","0101","0101","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","1000","0110","0110","0111","0111","0110","0110","0110","0101","0110","0101","0100","0100","0101","0111","0110","0101","0111","0111","0111","1000","1000","0110","0111","1000","1000","0110","0111","1000","1000","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0110","0111","0110","0110","0101","0100","0101","0101","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0100","0100","0110","0110","0100","0100","0011","0100","0100","0100","0100","0100","0011","0100","0101","0101","0011","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0101","0101","0101","0011","0001","0010","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0011","0100","0100","0011","0001","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0110","0100","0011","0100","0110","0110","0100","0101","0101","0101","0110","0101","0101","0011","0100","0100","0011","0011","0100","0100","0101","0100","0100","0100","0101","0101","0100","0011","0011","0100","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","1001","1001","1000","0110","0101","0110","1000","1001","1000","0110","1000","0111","0111","0110","1001","1001","1001","0110","0100","0101","1001","1001","1001","1001","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0110","0101","0101","0101","0101","0101","0101","0110","0111","0111","0111","1000","0110","0100","0100","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0101","0101","0111","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0101","0110","0110","0110","1000","0111","0111","1000","1000","0111","0111","1000","1000","0110","0111","1000","1000","0110","0101","0101","0101","0110","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0100","0100","0100","0101","0100","0101","0101","0101","0100","0101","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0011","0100","0100","0101","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0101","0011","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111"),
("0101","0101","0101","0010","0010","0001","0100","0101","0101","0110","0110","0110","0110","0101","0010","0010","0100","0110","0110","0101","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0100","0110","0111","0111","0110","0111","0111","0110","0110","0110","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","0101","0100","0011","0101","0110","0101","0101","0101","0101","0110","0110","0101","0100","0011","0100","0100","0011","0011","0100","0100","0100","0101","0100","0101","0101","0101","0101","0011","0011","0101","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","1000","1000","1000","0111","0110","0110","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1001","1001","1000","0101","0101","0110","1000","1000","1000","0110","0111","1000","0111","0110","1001","1001","1001","0110","0100","0101","1001","1001","1001","1001","1000","0110","0110","0111","1000","0111","0111","0111","1000","1000","0111","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","0111","0100","0100","0100","0101","0100","0100","0100","0100","0101","0111","0111","0111","0110","0100","0100","0100","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0101","0110","0110","0101","0101","0110","0101","0101","0101","0101","0101","0101","0100","0101","0101","0110","0111","0101","0101","0101","0100","0101","0111","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0110","0111","0111","1000","0111","0111","1000","1000","0111","0111","1000","1000","0111","0111","0111","1000","0110","0101","0101","0101","0101","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0110","0111","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0011","0101","1000","1000","0111","0111","0110","0111","1000","1000","1000","0111"),
("0110","0110","0101","0011","0010","0011","0100","0101","0101","0101","0101","0101","0110","0101","0010","0001","0011","0110","0110","0011","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0100","0010","0101","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0101","0011","0011","0101","0111","0110","0101","0101","0101","0110","0110","0101","0100","0011","0100","0100","0011","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0011","0011","0101","1011","1011","1010","1001","1001","1000","1000","1000","1000","1000","1000","1010","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","1000","0111","0111","0101","0101","0111","0111","0111","0111","0111","1000","1000","0111","0111","1000","1001","1001","1000","0101","0101","0110","1000","1001","1000","0110","0111","1000","0111","0110","1001","1010","1001","0110","0101","0101","1001","1001","1001","1001","0111","0110","0110","0111","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0111","0110","0110","0111","0111","0110","0100","0100","0100","0101","0101","0100","0100","0100","0101","0111","0111","0110","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0111","0111","0111","0111","0111","0101","0110","0110","0101","0101","0100","0101","0100","0100","0110","0111","0111","0100","0100","0101","0111","0111","0101","0100","0100","0110","0101","0110","1000","0111","0111","1000","1000","0111","0111","1000","1000","0110","0110","0101","0110","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0110","0101","0101","0100","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0110","1000","0110","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0011","0100","0111","0111","0111","0111","0101","0111","1000","1000","0111","0111"),
("0110","0110","0101","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0010","0001","0011","0110","0101","0011","0011","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0011","0110","0111","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","1000","1000","0111","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0101","0011","0011","0100","0110","0110","0110","0110","0101","0110","0101","0101","0100","0011","0100","0100","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0011","0011","0101","1010","1011","1010","1001","1001","1001","1000","1000","1000","1000","1001","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0110","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0110","0101","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1001","1001","1000","0101","0101","0110","1000","1000","1000","0110","1000","1000","0111","0110","1001","1010","1010","0110","0100","0101","1001","1001","1001","1001","1000","0110","0110","0110","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0110","0110","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0110","0101","0100","0101","0101","0101","0100","0100","0100","0101","0101","0100","0100","0100","0101","0110","0110","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0100","0101","0101","0100","0101","0101","0101","0101","0101","0110","0101","0110","0110","0110","0111","0111","0111","0101","0110","0101","0110","0110","0101","0101","0101","0101","0101","0100","0110","0110","0101","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0101","0111","1000","0111","0111","0111","1000","1000","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0111","0111","0111","0110","0111","0111","0111","0110","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0100","0101","0110","0101","0011","0100","0111","0111","0111","0111","0101","0100","0100","0100","0100","0011","0100","0011","0100","0011","0100","0100","0100","0100","0100","0110","0100","0100","1000","1000","0111","1000","0110","0111","1000","1000","1000","1000"),
("0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0010","0010","0011","0101","0110","0100","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0111","0111","0111","0111","0110","0100","0110","0111","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","0110","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0110","0100","0011","0100","0110","0110","0110","0110","0110","0110","0110","0101","0100","0011","0101","0101","0011","0100","0100","0101","0101","0101","0110","0110","0110","0110","0110","0011","0011","0101","1011","1011","1001","1001","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0110","0101","0110","0111","0111","1000","1000","0111","1000","1000","0111","0111","1000","1001","1001","1000","0101","0101","0110","1000","1001","1000","0110","0111","1000","0111","0110","1001","1010","1001","0110","0100","0110","1001","1001","1001","1001","0111","0101","0110","0101","0101","0111","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0111","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","0110","0110","0110","0110","0100","0100","0100","0100","0100","0100","0101","0110","0111","0111","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0111","0110","0110","0110","0110","0110","0110","0101","0101","0101","0110","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0101","0101","0101","0100","0100","0101","0100","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0111","0111","0111","0111","0111","0111","0110","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0101","0101","0100","0011","0011","0101","0101","0110","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0110","0101","0110","1000","1000","1000","1000","0111","0111","1000","1000","0111","0111"),
("0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0011","0010","0011","0101","0110","0100","0011","0101","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","1000","0111","0111","0111","0111","0111","0111","0110","1000","0111","0111","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0110","0100","0110","0110","0111","0111","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0111","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0100","0011","0101","0110","0110","0110","0110","0110","0110","0110","0101","0110","0101","0111","0111","0101","0101","0110","0101","0101","0110","0110","0110","0110","0110","0110","0100","0100","0110","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","1000","1001","1001","1000","0110","0101","0110","1000","1000","1000","0110","0111","1000","0111","0110","1001","1010","1010","0110","0100","0101","1001","1001","1001","1001","1000","0101","0110","0101","0100","0101","1000","1000","1000","1000","1000","0110","0111","0111","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0110","0110","0110","0110","0101","0110","0101","0101","0101","0110","0101","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0111","0111","0110","0111","0110","0111","1000","0111","0110","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0110","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0110","0110","0110","0110","0111","0110","0101","0101","0111","0111","0111","0110","0110","0110","0101","0101","0110","0101","0101","0111","0110","0101","0101","0110","0110","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0110","0101","0101","0101","0110","0110","0101","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0101","0110","0101","0101","0110","0110","0110","0110","0100","0101","0101","0101","0101","0100","0011","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0111","1000","1000","0101","0100"),
("0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0010","0001","0011","0101","0110","0100","0010","0101","0110","0110","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0110","0110","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0110","0110","0110","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0110","0011","0110","0111","0111","0110","0110","0110","0111","0110","0111","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","0111","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0111","0110","0111","1000","1001","1000","0111","0110","0100","0100","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0110","1000","0111","0110","0101","0111","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0101","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","0111","0111","1000","1000","0111","0111","1000","1000","1000","1000","1000","0110","0110","0110","0111","1000","0111","0111","1000","1000","1000","0111","0110","0101","0110","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0110","0101","0101","0111","0111","1000","1000","1000","1000","1000","0111","0111","1000","1001","1001","1000","0110","0101","0111","1000","1001","1000","0110","0111","1000","0111","0110","1001","1001","1010","0110","0100","0101","1001","1001","1001","1001","1000","0110","0111","0101","0100","0100","0111","0110","0111","0111","0111","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0110","0101","0101","0100","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0100","0111","1000","0111","0110","0110","1000","1000","0111","0110","0110","0110","0101","0101","0100","0101","0101","0100","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0100","0101","0110","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0100","0101","1000","0111","0110","0110","0111","0110","0101","0110","0111","0111","0111","1000","0100","0100","0110","0101","0100","0100","0110","0110","0101","0110","0111","0110","0110","0111","0110","0101","0100","0100","0100","0100","0100","0101","0101","0100","0101","0101","0110","0110","0101","0101","0101","0110","0110","0100","0100","0100","0100","0100","0101","0100","0100","0100","0101","0101","0100","0011","0011","0100","0100","0100","0100","0101","0100","0100","0101","0100","0100","0101","0101","0100","0011","0011","0011","0011","0100","0100","0011","0100","0101","0101","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0101","0100","0111","1000","1000","1000","1000","0111","1000","0111","0111","0101","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0101","0110","0101","0100","0011"),
("0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0010","0100","0101","0110","0100","0011","0101","0110","0110","0101","0101","0110","0110","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0111","1000","0111","0111","0111","0111","0111","0111","0110","0011","0101","0111","0111","0111","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0111","0111","0110","0110","0111","0111","0111","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","1000","0111","0110","0111","0110","0101","0110","0110","0110","0110","0101","0110","0110","0111","0111","1000","1001","1001","0111","0011","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0101","0110","0011","0011","0011","0011","0100","0110","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0100","0111","0111","0110","0110","0110","0110","0111","0111","0111","0110","0111","1000","0110","0110","0110","0110","0111","0111","1000","0111","1000","1000","1000","1000","1000","0111","0101","0110","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0110","0110","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0101","0101","0110","0111","0111","0111","0111","0111","0111","0110","0111","1000","1001","1001","1001","0110","0101","0110","1000","1000","1000","0110","0111","1000","0111","0110","1001","1010","1010","0110","0100","0101","1001","1001","1001","1001","1000","0110","0110","0101","0100","0100","0101","0110","0110","0110","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0110","0110","0110","0111","0110","0110","0110","0101","0110","0111","0111","0101","0101","0101","0101","0110","0110","1000","0111","1000","0111","0110","0111","0101","0110","0111","0101","0101","0110","0100","0100","0100","0101","0100","0111","1000","0111","0111","0111","1000","1000","0111","0110","0110","0101","0100","0100","0100","0100","0100","0101","0100","0101","0101","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0101","1000","1001","1000","0111","0110","0111","0110","0110","1000","1000","1000","1000","0101","0100","0110","0110","0100","0101","0111","0110","0101","0110","0111","0110","0111","0110","0110","0101","0100","0100","0100","0100","0100","0101","0101","0101","0100","0110","0110","0110","0101","0101","0101","0101","0110","0100","0011","0011","0011","0100","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0100","0100","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0011","0100","0101","0110","0101","0100","0100","0101","0100","0100","0101","0101","0101","0100","0100","0100","0101","0100","0100","0011","0011","0110","0111","1000","0111","1000","0110","0111","0111","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011"),
("0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0011","0001","0011","0101","0100","0011","0011","0100","0101","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0011","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","1000","1000","0111","0111","0111","0111","0110","0100","0011","0010","0011","0100","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0101","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0100","0100","0100","0100","0101","0110","0111","0110","0110","0110","0110","0111","0111","0111","0111","0101","0100","0100","0100","0100","0101","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","1000","1000","0111","1000","0111","0111","0111","1000","1000","0111","0111","1000","1000","0110","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0011","0101","0001","0001","0001","0001","0010","0101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0111","1000","1000","1000","1000","1000","1000","1000","0111","0111","0110","0110","0101","0110","0110","0110","0111","1000","1000","0111","1000","1000","0111","0110","0111","0110","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0110","0101","0101","0111","0111","1000","1000","1000","1000","1000","0111","0111","1000","1001","1001","1000","0110","0101","0110","1000","1000","1000","0110","0111","1000","0111","0110","1001","1010","1010","0111","0101","0101","1001","1001","1001","1001","1000","0110","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0101","0110","0111","0111","0110","0101","0110","0110","0101","0101","0101","0101","0101","1000","1010","0111","1001","1010","0111","0110","0110","0111","0111","0101","0110","0110","0100","0100","0100","0100","0100","0111","1000","0111","0110","0111","1000","1000","0111","0110","0101","0100","0100","0101","0101","0101","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0101","0111","0101","0111","1001","1000","0110","0101","0101","1000","0110","0110","1000","0101","0100","0101","0101","0100","0101","0111","0110","0101","0110","0111","0110","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0110","0110","1000","1000","0111","0101","0101","0100","0100","0011","0011","0100","0100","0101","0100","0011","0101","0101","0110","0110","0110","0101","0100","0011","0100","0100","0100","0100","0101","0100","0100","0101","0100","0100","0100","0100","0110","0111","0111","0111","0110","0100","0100","0101","0100","0101","0110","0101","0101","0101","0101","0100","0100","0110","0110","0100","0011","0011","0100","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0101","0101"),
("0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0011","0010","0100","0011","0010","0010","0010","0010","0011","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0100","0010","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0110","0110","0101","0011","0010","0010","0010","0010","0010","0011","0101","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0101","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0100","0100","0100","0100","0100","0110","0111","0110","0110","0110","0110","0111","0110","0110","0111","0101","0100","0100","0100","0101","0101","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","0111","0111","1000","0111","1000","0111","0111","0111","0101","0110","0110","0110","0110","0111","1000","1000","1000","0111","0110","1000","1001","0110","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0101","0010","0010","0010","0010","0011","0101","0010","0011","0011","0011","0011","0011","0011","0011","0011","0001","0001","0010","0110","0111","1000","1000","1000","0111","1000","1000","0111","1000","0111","0110","0101","0110","0110","0110","0111","1000","1000","0111","0111","1000","0110","0101","0111","0111","0101","0110","0111","0111","0111","0111","1000","1000","0111","0111","0110","0110","0110","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","1000","1001","1001","1000","0110","0101","0110","1001","1001","1000","0110","0110","0110","0111","0110","1001","1010","1001","0110","0100","0101","1001","1001","1001","1001","1000","0101","0110","0110","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1001","0111","1000","1001","0111","0101","0101","0101","0111","0101","0110","0110","0111","1010","0111","1001","1001","0110","0111","0110","0111","1000","0110","0111","0110","0100","0101","0100","0100","0100","0111","1000","0111","0110","0111","0111","1000","0111","0101","0101","0101","0100","0101","0101","0101","0101","0101","0110","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","1000","1000","1001","1010","1001","0111","0101","0101","1000","1000","1001","1000","0101","0101","0101","0101","0100","0101","0111","0110","0101","0110","0110","0110","0110","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0101","0101","0111","1000","0111","0101","0100","0100","0101","0011","0100","0100","0101","0110","0101","0011","0100","0101","0101","0110","0101","0011","0011","0011","0011","0100","0011","0100","0100","0011","0011","0101","0100","0100","0101","0110","0111","0110","0110","0110","0110","0101","0011","0101","0101","0110","0101","0101","0101","0101","0101","0011","0100","0100","0100","0011","0011","0011","0011","0100","0101","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0011","0011","0100","0101","0101","0101","0100"),
("0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","1000","0111","0110","0110","0110","0011","0010","0010","0010","0010","0010","0010","0010","0011","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0111","0111","0111","0111","0110","0111","0111","0110","0110","0110","0110","0110","0101","0101","0101","0101","0110","0101","0100","0110","0101","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0111","0111","0111","0111","0110","0111","0110","0110","0111","0111","0111","0111","0111","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0100","0101","0110","0110","0101","0101","0101","0110","0101","0110","0110","0110","0110","0110","0111","1001","1001","1001","1000","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","0111","0111","0110","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","1000","1001","0110","0010","0010","0011","0101","0101","0101","0100","0101","0101","0101","0100","0100","0101","0010","0011","0011","0010","0011","0101","0100","0100","0101","0101","0100","0100","0101","0101","0100","0010","0010","0011","0110","1000","1001","1001","1001","1001","1001","1001","1000","1000","0111","0110","0110","0110","0110","0111","1000","1000","1000","1000","1000","1000","0110","0100","0101","0101","0101","0101","0111","0111","0111","0111","1000","1000","0111","0111","0110","0110","0110","0110","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0110","0110","0111","0111","1000","1000","1000","0111","0111","0111","0110","1000","1001","1001","1001","0110","0100","0110","1000","1001","1000","0110","0110","0101","0101","0110","0111","0111","1000","0110","0101","0101","1001","1010","1001","1001","1000","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1001","1000","1001","1010","0110","0110","0110","0110","0111","0110","0110","0110","1000","1010","0111","1001","1010","0110","0101","0101","0110","0111","0110","0111","0110","0100","0100","0100","0100","0101","0110","0111","0110","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0100","0100","0101","0101","0100","0100","0101","0110","0111","0110","0110","0101","0101","0101","0110","0101","0100","0100","0100","0101","0100","0100","0100","1000","1001","1001","1010","1001","1000","1000","1000","1000","1000","1000","0111","0101","0101","0101","0100","0100","0101","0110","0101","0101","0101","0110","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0100","0100","0101","0110","0110","0111","0111","0111","0111","0110","0100","0100","0100","0101","0101","0101","0110","0110","0110","0101","0011","0100","0101","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0101","0110","0101","0101","0100","0100","0101","0110","0101","0100","0101","0101","0100","0100","0100","0100","0100","0101","0011","0100","0100","0100","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0100","0110","0101","0101","0100","0101","0100","0100","0011","0011","0100","0100","0100","0100","0011","0011"),
("0101","0101","0101","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","1000","1000","0111","0110","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0100","0100","0101","0100","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0110","0110","0110","0101","0101","0101","0101","0101","0110","0110","0110","0101","0110","0110","0110","0101","0101","0101","0101","0101","0110","0110","0101","0110","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0101","0110","0101","0101","0100","0100","0011","0100","0101","0110","0110","0111","0111","0111","0111","0101","0110","0110","0110","0111","1000","1001","1001","1001","1001","1000","1000","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0110","0111","0110","0110","0110","0110","0111","0111","1000","1000","0111","1000","1000","0101","0010","0010","0100","0110","0101","0100","0010","0100","0101","0101","0100","0101","0110","0011","0011","0100","0011","0100","0101","0011","0100","0101","0101","0011","0011","0100","0101","0101","0011","0010","0011","0101","1000","1000","1000","1000","1000","1001","1000","1000","1000","0111","0110","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0110","0100","0100","0101","0101","0101","0111","0111","1000","0111","1000","1000","1000","0111","0101","0101","0110","0110","0111","0110","0111","0111","0111","1000","0111","0111","0111","0111","0111","0101","0101","0111","0111","1000","0111","0111","0101","0110","0110","0110","0111","0111","1000","1000","0101","0100","0100","0111","1000","0111","0110","0110","0101","0101","0110","0111","0111","0110","0110","0101","0101","1000","1001","1001","1000","0110","0101","0110","0110","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1000","0111","0111","1000","0110","0111","1000","0111","1000","0110","0111","0111","0110","0111","0110","1001","1010","0111","0111","0110","0110","0110","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0110","0110","0101","0100","0100","0101","0101","0100","0100","0110","0101","0101","0100","0100","0100","0101","0111","0110","0100","0100","0100","0011","0100","0100","0100","1000","1000","1001","1000","1000","1001","1001","1001","1001","1001","1001","1000","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0101","0110","0111","0111","0111","0101","0101","0101","0100","0011","0100","0101","0110","1000","0111","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0011","0100","0100","0100","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0101","0110","0101","0101","0011","0100","0100","0100","0100","0011","0100","0101","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0100","0100","0100","0100","0101","0011","0011","0100","0100","0100","0100","0011","0011"),
("0101","0101","0101","0101","0100","0100","0100","0101","0100","0101","0101","0101","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0111","1000","1000","0111","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0111","0110","0111","0111","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0111","0110","0111","0110","0111","0111","0111","0110","0101","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0101","0101","0110","0111","0110","0100","0101","0101","0110","0111","0110","0101","0101","0101","0111","0110","0101","0101","0101","0110","0111","0111","0110","0110","0110","0111","0111","1000","0111","0111","0111","1000","0111","1000","0111","0111","1000","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0110","0110","0101","0100","0100","0100","0101","0101","0110","0110","0101","0100","0100","0100","0100","0101","0110","0110","0110","0110","0110","0110","0101","0110","0111","0111","0110","1000","1001","1001","1001","1001","1000","1000","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","1000","1000","0101","0011","0011","0100","0110","0101","0101","0010","0100","0101","0101","0100","0101","0110","0011","0100","0100","0011","0101","0101","0100","0100","0101","0101","0011","0011","0101","0101","0101","0011","0010","0011","0101","1000","1000","1000","1000","0111","1001","1000","1000","0111","0111","0110","0101","0101","0110","0101","0111","1000","1000","1000","1000","0110","0100","0100","0100","0101","0101","0101","0111","0111","0111","0111","0111","0111","0111","0110","0101","0101","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0100","0101","0111","0111","0111","0110","0101","0100","0101","0101","0101","0101","0101","0110","0101","0100","0100","0101","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","1001","0111","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0110","1000","0111","0110","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0100","0101","0100","0011","0011","0100","0101","0110","0110","0101","0101","0110","0110","0110","0101","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0110","0101","0101","0100","0100","0100","0100","0100","0100","0101","1000","0111","1000","1000","0110","0101","0110","1001","0111","0101","0111","0111","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0111","0110","0111","0101","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0011","0011","0100","0100","0101","0101","0100","0101","0101","0101","0101","0100","0100","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011"),
("0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0101","0110","0110","0101","0110","0101","0101","0101","0101","0110","0110","0110","0110","0111","0110","0111","0111","0111","0111","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0101","0101","0110","0110","0110","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0101","0110","0111","0111","0111","1000","1000","0111","0111","0111","0111","1000","0111","0111","1000","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0110","0110","0100","0100","0100","0101","0101","0110","0110","0110","0101","0100","0100","0100","0101","0110","0110","0101","0100","0100","0101","0110","0110","0110","0111","0111","0111","1000","1001","1001","1001","1001","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","0110","0111","0110","0110","0110","0110","0110","0110","0111","0111","1000","0111","0110","1000","1000","0101","0011","0011","0101","0111","0110","0110","0100","0101","0110","0111","0101","0110","0110","0100","0100","0100","0100","0110","0110","0101","0100","0101","0101","0011","0100","0110","0101","0101","0011","0010","0100","0101","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0110","0101","0110","0101","1000","1000","1000","0111","0111","0110","0100","0100","0100","0101","0101","0101","0111","0111","0111","1000","1000","1000","0111","0101","0100","0101","0110","0110","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0100","0101","0101","0101","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0100","0100","0100","0101","0110","0111","0111","0110","0110","0110","0101","0101","0110","0110","0111","0110","0111","0110","0100","0100","0100","0100","0100","0101","0101","0101","0111","0111","0111","0111","0110","0110","0100","0011","0011","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0101","0101","0100","0100","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0101","0111","1000","0101","0101","0100","0011","0011","0011","0101","0101","0101","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0101","0100","0100","0110","0101","0101","0110","0101","0101","0110","1000","0110","0110","0110","0110","0101","0101","0111","0101","0100","0101","0110","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0110","0110","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0101","0100","0011","0011","0011","0011","0011"),
("0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0111","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0111","0111","0111","0110","0101","0110","0111","0111","0110","0100","0101","0110","0111","0111","0101","0101","0110","0111","0111","0111","0101","0110","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0100","0100","0101","0111","0110","0110","0111","0111","0110","0100","0100","0100","0100","0110","0110","0101","0100","0100","0101","0101","0101","0110","0111","0111","0110","1000","1001","1001","1001","1001","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1001","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","1000","1000","1000","0111","0101","0111","0110","0100","0011","0011","0100","0110","0110","0111","0100","0100","0111","0111","0101","0101","0100","0011","0100","0101","0100","0100","0100","0100","0101","0101","0101","0100","0101","0110","0110","0110","0011","0010","0011","0011","0101","1000","1000","0111","0111","1000","1000","1000","1000","0111","0110","0110","0110","0110","0110","1000","1000","1000","0110","0111","0101","0100","0100","0100","0100","0100","0101","0110","0110","0110","0111","0110","0110","0101","0101","0100","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0101","0110","0110","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0110","0101","0101","0100","0101","0100","0100","0100","0100","0110","0101","0111","1000","1000","0110","0100","0110","1000","1000","1000","1000","0111","0110","0110","0101","0101","0111","0111","0111","0110","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0101","0100","0101","0101","0101","0100","0110","0110","0100","0101","0100","0100","0100","0100","0111","0111","0111","0101","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0101","0110","0110","0110","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0110","0110","0101","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0011","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011"),
("0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0001","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0100","0101","0101","0101","0101","0101","0100","0101","0100","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0011","0011","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0111","0110","0111","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0110","0110","0110","0110","0110","0111","0110","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0101","0110","0110","0101","0101","0100","0101","0110","0101","0101","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0101","0110","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0110","0110","0100","0100","0100","0100","0101","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0101","0100","0101","0101","0101","0110","0110","0110","0111","0110","1000","1001","1001","1001","1001","1000","0111","0111","0111","0111","0111","1000","0111","0111","0111","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0110","1000","1000","0111","0111","0111","0111","1000","0110","0100","0110","0100","0011","0010","0010","0100","0111","0101","0101","0101","0101","0110","0111","0101","0100","0100","0011","0100","0101","0100","0100","0100","0100","0101","0110","0110","0101","0101","0011","0101","0110","0010","0001","0011","0100","0110","1000","1000","1000","1000","1001","1000","1000","1000","0111","0100","0101","0110","0110","0101","0110","0101","0111","0110","0101","0100","0100","0100","0100","0100","0101","0110","0110","0101","0101","0110","0110","0110","0110","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0100","0101","0101","0100","0111","1000","0111","0111","0111","0110","0110","0111","0111","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","0110","0111","0111","0111","0111","1000","0111","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0011","0010","0101","1010","1010","1010","1010","1001","1000","0111","0110","0101","0110","0111","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0110","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0110","0101","0100","0100","0101","0111","0110","0111","0110","0101","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0110","0111","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0100","0101","0101","0110","0101","0110","0110","0101","0110","0110","0101","0101","0100","0101","0111","1000","1000","0101","0100","0101","0101","0100","0100","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0011","0101","0101","0100","0011","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0011","0011","0011"),
("0100","0100","0100","0100","0100","0100","0101","0100","0101","0101","0101","0101","0101","0100","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0100","0100","0101","0110","0111","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0110","0011","0001","0010","0001","0010","0010","0011","0010","0010","0010","0011","0001","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0101","0110","0110","0101","0110","0110","0110","0110","0101","0101","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0110","0111","0111","0111","0111","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","1000","0110","0110","0101","0110","0111","0111","0110","0101","0101","0111","0111","0111","0101","0101","0101","0111","0111","0110","0110","0110","0111","0111","0111","0101","0110","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0101","0100","0100","0011","0100","0110","0111","0111","0110","0100","0100","0100","0100","0110","0110","0101","0100","0100","0100","0100","0101","0111","0111","0111","0110","0111","1001","1001","1001","1001","1000","0111","0111","0101","0101","0111","1000","1000","0111","0111","1000","1000","0111","0110","0110","0110","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","1000","1000","0101","0100","0100","0101","0100","0010","0010","0100","0110","0011","0100","0101","0101","0110","0110","0100","0101","0101","0011","0101","0110","0100","0100","0101","0100","0101","0110","0110","0101","0101","0011","0100","0110","0011","0010","0011","0100","0101","0110","0110","0110","0110","1000","0111","0111","0111","0110","0101","0101","0110","0111","0111","0101","0100","0110","0110","0100","0100","0100","0100","0100","0100","0101","0110","0110","0101","0101","0110","0110","0111","0111","0110","0100","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0110","0110","0110","0101","0100","0100","0101","0101","0101","0100","0100","0101","0101","0111","0111","0111","0111","1000","0111","0110","0101","0101","0110","0101","0101","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","1000","1001","1001","1001","0111","0111","0111","0110","0101","0110","0110","0101","0101","0101","0100","0101","0101","0100","0100","0100","0110","0101","0101","0101","0110","0101","0101","0111","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0101","1001","1001","0111","0110","0100","0011","0011","0011","0011","0011","0100","0100","0101","0101","0101","0110","0110","0111","0111","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0101","0101","0101","0101","0100","0011","0100","0100","0101","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0010","0010","0010","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0110","0110","0101","0100","0101","0110","1000","0111","0111","0110","0110","0111","0110","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","1000","1000","1000","1000","0111","0110","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0011","0011"),
("0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0010","0010","0010","0010","0001","0100","0100","0001","0001","0010","0011","0001","0011","0100","0101","0110","0110","0110","0110","0110","0101","0100","0100","0100","0100","0011","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0100","0010","0100","0010","0001","0011","0110","0011","0001","0010","0100","0010","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0110","0110","0110","0101","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0101","0101","0101","0110","0110","0110","0101","0101","0110","0111","0111","0110","0101","0100","0101","0110","0111","0101","0101","0101","0110","0110","0110","0101","0110","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0110","0110","0110","0111","0111","0101","0101","0110","0110","0110","0110","0101","0100","0101","0101","0101","0110","0101","0101","0100","0101","0101","0110","0110","0110","0110","0110","0111","1001","1001","1001","1001","0111","0110","0101","0100","0100","0101","0111","0111","0110","0110","0110","0110","0110","0101","0100","0100","0110","1000","0111","0111","0110","0110","0101","0101","0110","0101","0101","0110","0111","0101","0100","0100","0101","0100","0010","0010","0100","0101","0011","0011","0101","0101","0110","0110","0101","0101","0101","0100","0101","0111","0101","0101","0101","0100","0101","0110","0101","0101","0100","0011","0011","0101","0011","0010","0011","0100","0100","0110","0111","0110","0101","0111","0110","0111","0110","0110","0111","0111","0111","0111","1000","0101","0100","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0101","0110","0101","0110","0110","0101","0110","0101","0101","0101","0100","0100","0101","0111","0111","1000","0111","0111","0110","0111","0110","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0110","0110","0110","0111","0101","0110","0101","0100","0100","0101","0101","0101","0100","0100","0100","0100","0101","0110","0110","0111","1000","1000","0101","0100","0100","0101","0101","0100","0011","0011","0100","0101","0100","0100","0100","0100","0110","0111","0111","0100","0100","1000","1001","1001","1001","0111","0110","0111","0101","0100","0110","0111","0101","0101","0101","0100","0100","0100","0100","0100","0100","0110","0100","0101","0101","0110","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0111","0101","0101","0100","0011","0011","0100","0011","0011","0011","0100","0100","0110","0110","0101","0101","0101","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0101","0100","0100","0100","0100","0100","0100","0100","0101","0011","0011","0010","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0010","0011","0110","0110","0101","0101","0101","0110","0100","0101","0111","0101","0110","0100","0011","0100","0101","0100","0101","0100","0101","0100","0110","0111","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0101","0101","0100","0101","0101","0100","0100","0100","0100","0011","0011","0100","0011","0100","0011","0011","0011","0100","0110","0110","0110","0111","0111","0101","0100","0100","0100","0101","0100","0100","0101","0101","0100","0100","0100","0100","0101","0101","0100","0100","0101","0100","0011","0011","0100","0101","0110","0101","0110","0101","0011","0101","0100","0100","0101","0100","0100","0100","0101","0011","0011","0011","0011"),
("0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0010","0010","0010","0010","0001","0010","0011","0001","0001","0010","0010","0010","0011","0100","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0100","0101","0100","0100","0100","0100","0101","0101","0100","0100","0101","0110","0100","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0111","0110","0110","0110","0110","0111","0111","0111","0111","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0101","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0101","0101","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0110","0110","0110","0101","0110","0101","0110","0111","1000","1000","0111","0101","0100","0101","0111","0111","0110","0110","0110","0111","0111","0111","0101","0110","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0101","0100","0100","0100","0100","0110","0110","0101","0100","0100","0101","0111","0110","0111","0111","0111","0111","1000","1001","1001","1001","1000","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0011","0100","0111","0111","0111","0111","0111","0111","0111","0111","0101","0100","0110","0110","0100","0100","0100","0101","0100","0011","0010","0100","0100","0011","0101","0101","0101","0101","0111","0101","0100","0101","0100","0101","0111","0100","0100","0100","0100","0101","0110","0110","0110","0101","0101","0011","0011","0011","0011","0011","0100","0101","1000","1000","1000","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","1000","1000","1000","0110","0110","0110","0110","0110","0110","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0111","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","0111","0110","0100","0011","0100","0100","0100","0100","0100","0101","0100","0110","0101","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0110","0110","1000","1000","0111","0101","0100","0100","0101","0101","0100","0100","0011","0100","0101","0101","0100","0100","0101","1001","1000","1001","0110","0101","1000","1001","1001","1001","0111","0110","0110","0100","0011","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0110","0100","0100","0110","0101","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0110","0101","0101","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0010","0010","0110","0111","0110","0110","0110","1000","0110","0110","0110","0101","0110","0100","0010","0100","0110","0101","0110","0101","0110","0101","0111","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0100","0101","0101","0101","0110","1000","0110","0101","0101","0101","0110","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0101","0100","0100","0101","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0010","0011","0010","0011","0011","0011","0011","0011","0011","0100","0110","0110","0110","0110","0110","0110","0110","0011","0011","0011","0011"),
("0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0010","0001","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0011","0100","0101","0101","0101","0101","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0100","0100","0100","0100","0101","0100","0100","0101","0110","0100","0001","0010","0010","0010","0010","0011","0010","0010","0010","0010","0001","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0101","0101","0110","0110","0101","0100","0100","0101","0101","0101","0101","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0101","0110","0110","0110","0110","0110","0101","0101","0110","0110","0110","0111","1001","1000","0110","0110","0101","0100","0100","0101","0111","0111","0111","0110","0110","0110","0110","0111","1000","1000","0111","0111","0111","0111","0110","0111","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0111","1000","1000","0110","0101","0100","0101","0101","0111","0110","0110","0101","0110","0110","0111","0101","0110","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0111","0110","0110","0111","0111","0110","0110","0111","0111","0110","0110","0101","0100","0100","0101","0110","0110","0110","0101","0101","0101","0100","0100","0100","0110","0110","0101","0101","0101","0101","0110","0110","0111","0111","0111","0111","1000","1001","1001","1001","1000","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0011","0100","0110","0101","0101","0101","0110","0111","0111","0111","0101","0100","0101","0101","0100","0100","0100","0101","0100","0011","0010","0100","0011","0100","0011","0101","0101","0101","0101","0100","0100","0100","0011","0100","0110","0100","0100","0100","0100","0100","0101","0101","0110","0011","0010","0100","0011","0011","0011","0011","0100","0110","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1001","1000","1001","1000","1001","1000","1000","1000","1001","1001","1001","1000","0110","0110","0110","0110","0111","0110","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0111","1000","1000","0110","0110","0110","1000","0111","0110","0111","1000","1001","0110","0100","0110","0101","0100","0011","0100","0101","0100","0100","0101","0111","0110","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0110","0110","0110","0111","0111","0110","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0101","1000","0101","0111","0101","0100","1000","1001","1001","1001","0111","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0110","0110","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0010","0010","0010","0100","0101","0101","0101","0101","0101","0101","0110","0110","0101","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0010","0010","0010","0101","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0100","0011","0100","0111","0111","0111","0111","0111","0110","0110","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0100","0100","0100","0100","0101","0100","0010","0011","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0110","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0110","0110","0110","0101","0110","1000","0110","0011","0011","0011","0011"),
("0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0010","0010","0010","0010","0001","0011","0100","0001","0001","0010","0010","0001","0011","0100","0101","0101","0101","0101","0100","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0101","0101","0100","0100","0101","0110","0100","0010","0100","0010","0001","0011","0110","0011","0001","0010","0100","0010","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0101","0110","0110","0110","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0111","0111","0110","0111","1000","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0100","0110","0110","0101","0101","0100","0101","0101","0101","0100","0101","0100","0110","0111","1000","1000","0111","0111","0111","0110","0101","0101","0111","0111","0110","0110","0101","0101","0110","0111","0111","0111","0111","0111","0111","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0011","0100","0110","0111","0110","1000","1001","1000","0111","0101","0101","0101","0111","0111","0110","0101","0101","0110","0111","0111","0110","0110","0111","0111","1000","1000","0111","0111","0110","0110","1000","0111","0101","0110","0101","0100","0110","1000","0111","1000","0111","0110","0110","1001","0111","0111","0110","0101","0100","0100","0100","0100","0110","0111","0110","0101","0100","0100","0100","0101","0110","0110","0101","0100","0100","0100","0100","0110","0111","0111","0111","0111","1000","1001","1001","1001","1000","0100","0101","0101","0100","0101","0111","0111","0110","0110","0101","0100","0101","0101","0101","0101","0011","0011","0100","0101","0110","0110","0110","0110","0111","0110","0100","0100","0100","0101","0100","0100","0110","0101","0100","0011","0010","0011","0100","0011","0001","0010","0101","0110","0101","0100","0100","0101","0100","0100","0110","0011","0100","0100","0100","0100","0100","0100","0011","0001","0001","0010","0011","0011","0011","0011","0100","0101","0110","0110","0110","0110","0110","1000","1000","1000","1001","1000","1001","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","0111","0111","0110","0111","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0111","1000","0111","0110","0110","0101","0110","0110","0101","0111","1000","1000","0110","0101","0101","0101","0100","0011","0100","0101","0101","0101","0101","0110","0111","0110","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0110","0111","0111","0100","0011","0011","0011","0011","0011","0011","0100","0100","0101","0110","1000","0101","1000","0110","0100","1000","1000","1001","1001","0111","0100","0100","0101","0101","0100","0100","0100","0100","0100","0011","0100","0101","0101","0101","0101","0011","0011","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0101","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0101","0100","0011","0100","0100","0100","0100","0100","0100","0110","0100","0100","0100","0100","0100","0011","0011","0011","0100","0101","0110","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0011","0010","0011","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0110","0101","0101","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0100","0100","0100","0101","0110","0100","0010","0101","0111","0100","0110","0101","0101","0101","0110","0101","0111","1000","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0111","0111","0110","0111","0111","1000","0110","0100","0011","0011","0011"),
("0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0010","0011","0010","0001","0011","0100","0010","0001","0010","0010","0010","0011","0100","0101","0101","0101","0101","0101","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0101","0100","0100","0101","0110","0100","0010","0100","0010","0001","0011","0110","0100","0001","0010","0100","0010","0011","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0101","0100","0100","0101","0110","0110","0110","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","0110","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0110","0110","1000","1000","1001","1001","1000","0110","0111","1001","1001","1001","1001","0111","0101","0101","0100","0011","0101","0100","0101","0101","0101","0101","0110","1000","0110","0100","0110","0111","0111","0110","0101","0100","0100","0100","0100","0100","0100","0100","0101","0111","1000","1000","0111","0111","1000","1000","0111","0110","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","1000","0111","0110","0100","0101","1000","0110","0110","0101","0100","0100","0111","1001","1001","1000","0111","1000","1001","1000","1000","0110","0101","0100","0100","0100","0101","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0101","0101","0100","0101","0110","0111","0111","0111","0110","0111","1001","1001","1001","1000","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0100","0110","0110","0110","0111","0111","0111","0101","0100","0100","0100","0100","0100","0100","0101","0110","0101","0011","0011","0011","0011","0010","0001","0000","0100","0110","0101","0101","0101","0101","0100","0100","0101","0100","0100","0101","0101","0101","0101","0101","0010","0000","0001","0001","0011","0011","0011","0011","0101","0101","0101","0101","0101","0101","0100","0101","0110","0110","0110","0110","0111","0110","0110","0110","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0110","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0110","0111","0110","0110","0110","0101","0101","0100","0110","0111","0101","0101","0101","0110","0111","0111","0111","0101","0101","0101","0100","0101","0100","0100","0101","0101","0101","0100","0100","0110","0110","0110","0110","0101","0101","0100","0011","0011","0011","0011","0100","0101","0101","0110","1001","0101","1000","0110","0101","1001","1000","1000","1010","1000","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0011","0011","0100","0101","0101","0110","0101","0100","0100","0100","0100","0100","0100","0100","0101","0110","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0101","0101","0100","0011","0100","0100","0100","0100","0100","0100","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0100","0110","0110","0101","0100","0100","0100","0100","0011","0011","0100","0101","0100","0011","0100","0100","0100","0100","0011","0100","0011","0100","0100","0100","0011","0011","0011","0011","0101","0110","0101","0011","0010","0100","0101","0101","0110","0101","0101","0110","0110","0110","1000","0110","0101","0101","0100","0101","0110","0111","1000","0111","0100","0101","0101","0100","0100","0100","0101","0110","0110","0110","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0111","0111","0111","0110","0110","0110","0110","0100","0011","0011","0010"),
("0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0010","0010","0011","0010","0001","0011","0100","0010","0001","0010","0011","0001","0011","0100","0101","0101","0101","0101","0101","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0011","0011","0100","0100","0100","0101","0110","0100","0010","0100","0010","0001","0010","0110","0100","0001","0010","0100","0010","0011","0110","0111","0111","0110","0110","0110","0110","0101","0101","0101","0101","0100","0100","0101","0110","0110","0111","0110","0101","0110","0110","0110","0110","0110","0111","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0110","0110","0110","0101","0100","0011","0010","0100","0100","0011","0011","0011","0100","0100","0101","0110","1000","1001","1001","1001","1001","1001","1001","1001","1010","0111","0100","0100","0011","0011","0101","0100","0100","0100","0101","0101","0101","0101","0100","0011","0100","0101","0110","0110","0101","0100","0100","0100","0100","0100","0101","1000","1001","1011","1011","1011","1010","1001","1000","1000","1000","0111","0101","0110","0110","0111","1000","0111","0101","0101","0110","0111","0111","0110","0110","0111","1000","0111","0111","0110","0101","0100","0101","0110","0100","0101","0100","0100","0100","0111","1001","1001","0111","0100","0101","1000","1000","1000","0110","0110","0100","0100","0101","0110","0110","0110","0111","0110","0110","0111","0111","0111","0111","0110","0110","0101","0100","0100","0101","0110","0110","0111","0110","0111","0110","0111","1001","1001","1001","1000","0101","0101","0100","0011","0101","0111","0110","0111","1000","0111","0111","1000","0111","0110","0100","0100","0011","0100","0110","0111","0110","0111","0111","0111","0101","0100","0011","0100","0100","0100","0100","0101","0111","0110","0100","0011","0011","0011","0010","0001","0001","0011","0110","0101","0110","0111","0111","0101","0101","0101","0100","0101","0111","0110","0101","0110","0101","0010","0000","0001","0010","0010","0011","0011","0100","0111","0111","0101","0101","0100","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0110","0111","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","0111","0110","0110","0101","0100","0100","0100","0100","0100","0100","0110","0100","0100","0100","0100","0101","0100","0100","0011","0011","0100","0110","0101","0101","0101","0101","0110","0101","0100","0100","0100","0101","0110","0110","0110","0101","0101","0100","0101","0101","0110","0100","0101","0101","0101","0101","0101","0100","0101","0100","0100","0101","0101","0110","0110","0110","0101","0101","0101","0011","0011","0011","0011","0011","0101","1000","1000","1010","1001","1010","0110","0101","0110","0100","0100","0111","0110","0101","0111","1000","0110","0101","0101","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0011","0011","0100","0100","0110","0111","0101","0011","0011","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0100","0011","0011","0100","0100","0011","0100","0110","0110","1000","1001","0110","0100","0011","0100","0100","0011","0011","0101","0101","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0110","0110","0110","0110","1000","1000","1000","1000","0110","0101","0101","0101","0101","0101","0101","0110","0101","0100","0011","0011","0010","0011","0011","0100","0101","0100","0100","0100","0100","0100","0100","0011","0100","0101","0100","0010","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0100","0100","0011","0010","0010","0001","0100","1001","1000","0101","0101","0101","0110","1001","0110","0101","0101","0101","0101","0101","0100","0110","0110","0110","0100","0100","0100","0100","0100","0100","0110","0110","0110","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0110","0110","0111","0100","0011","0100","0101","0011","0011","0011","0010"),
("0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0010","0010","0011","0010","0001","0011","0100","0010","0001","0010","0010","0001","0011","0100","0101","0101","0101","0101","0101","0100","0011","0011","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0011","0100","0100","0100","0100","0100","0100","0100","0101","0110","0100","0010","0100","0010","0001","0010","0101","0100","0010","0001","0100","0010","0011","1000","1000","0111","0111","0111","0110","0110","0110","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0101","0101","0110","0110","0110","0101","0110","0101","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","1000","1000","1000","1000","0111","0110","0011","0010","0101","0101","0011","0100","0101","0100","0100","0100","0101","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0100","0011","0011","0100","0110","0110","0111","0110","0110","0110","0110","0111","0101","0011","0100","0101","0101","0101","0101","0100","0100","0100","0100","0101","1001","1010","1011","1010","1001","1001","1010","1010","1001","1001","1000","0111","1000","0111","1000","0111","1001","0111","0101","0110","0110","0111","0111","0110","0110","0111","1000","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0111","1010","1001","0111","0101","0101","0101","1001","1000","0110","0101","0110","0111","0111","0111","0110","0110","0110","0110","0110","0111","0111","0111","0110","0101","0101","0100","0011","0100","0100","0101","0101","0101","0110","0110","0110","1000","1001","1001","1001","1000","0101","0100","0100","0011","0101","0111","0111","1000","1000","0111","0111","0111","0111","0101","0100","0100","0100","0100","0101","0111","0110","0110","0101","0101","0101","0110","0100","0011","0011","0011","0101","1000","1010","0111","0101","0011","0011","0010","0010","0001","0010","0010","0100","0101","0111","1001","1001","0111","0110","0111","0110","0110","1000","1000","0110","0101","0011","0001","0001","0001","0010","0010","0100","0011","0100","0111","1001","0111","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0100","0011","0100","0101","0100","0101","0101","0110","0101","0101","0110","0110","0110","0110","0111","0111","0101","0101","0110","0101","0100","0100","0100","0101","0100","0100","0011","0101","0101","0101","0110","1000","0100","0011","0011","0011","0100","0101","0101","0101","0101","0100","0100","0011","0011","0100","0101","0111","1001","0101","0100","0100","0100","0100","0100","0100","0101","0100","0110","0111","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0111","0110","0101","0011","0011","0011","0011","0100","0101","0111","0111","1010","1001","1011","0111","0011","0011","0100","0100","0100","0100","0100","0110","1001","0110","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0101","0100","0011","0011","0100","0110","0110","0110","0110","0110","0110","0110","0101","0101","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0110","0111","0111","0100","0100","0101","0101","0110","1000","0111","0101","0100","0100","0100","0100","0100","0100","0110","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0100","0011","0011","0100","0111","1000","1000","1000","0110","0100","0100","0101","0101","0101","0100","0101","0100","0100","0011","0010","0010","0010","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0101","0101","0100","0100","0100","0111","0111","0101","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0110","0110","0101","0101","0101","0100","0101","0011","0011","0101","0110","0101","0101","0110","0101","0100","0010","0011","0101","0101","0011","0011","0101","0100","0011","0110","0110","0101","0100","0100","0100","0011","0011","0011","0010","0010"),
("0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0101","0101","0100","0010","0010","0100","0010","0010","0010","0100","0010","0001","0010","0011","0001","0011","0100","0101","0101","0101","0101","0101","0100","0100","0100","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0010","0100","0010","0001","0010","0100","0101","0011","0001","0100","0010","0011","0111","0111","0110","0110","0111","0110","0101","0110","0101","0101","0101","0110","0101","0101","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0110","0110","0110","0110","0111","0110","0100","0101","0110","0101","0101","0110","0101","0110","0111","0101","0101","0101","0101","0101","0011","0100","0101","0101","0011","0011","0100","0100","0100","0100","0100","0111","0110","0101","0110","1001","1010","1001","1001","1001","1001","0111","0011","0011","0011","0101","0101","0101","0101","0101","0110","0111","0111","0110","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0101","0110","0110","0110","0111","1001","1010","1001","1001","1000","0111","1001","0110","1000","0111","1010","0111","0101","0101","0110","0110","0110","0110","0110","0111","1000","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0111","1001","1001","0111","0100","0100","0101","1000","1000","0111","0110","0110","0111","0110","0111","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0100","0100","0101","0101","0101","0110","0110","0110","0111","1000","1000","0110","0100","0100","0100","0100","0100","0100","0110","1000","1000","0110","0101","0101","0110","0101","0100","0011","0100","0100","0101","0111","0110","0110","0101","0101","0110","1000","0110","0101","0101","0110","0111","0111","0110","0100","0011","0011","0100","0010","0010","0001","0011","0011","0100","0100","0101","0101","0100","0100","0100","0101","0011","0100","0100","0100","0100","0100","0011","0001","0001","0001","0010","0010","0101","0100","0010","0010","0011","0100","0101","0101","0101","0110","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0110","0110","0111","0101","0101","0100","0100","0100","0011","0011","0010","0011","0100","0101","0101","0111","1001","0011","0011","0011","0011","0011","0100","0110","0110","0101","0101","0101","0100","0100","0100","0100","0110","1010","0100","0011","0011","0011","0100","0100","0100","0101","0100","0110","0110","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0110","0101","0011","0100","0100","0100","0100","0101","0110","0110","1001","0111","1001","1001","0111","0111","0111","0111","0111","0111","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0011","0100","0100","0101","0110","0111","0011","0001","0001","0001","0011","0110","0101","0100","0100","0100","0100","0100","0100","0100","0101","0110","0110","0110","0111","0111","1000","0110","0100","0101","1000","0111","0101","0101","0101","0101","0101","0101","0101","0101","0111","1000","0101","0011","0110","1000","0011","0010","0010","0011","0100","0100","0100","0110","0101","0100","0110","0110","0101","0101","0100","0100","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0101","0101","0101","0101","0101","0100","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0001","0010","0100","0100","0100","0011","0011","0100","0100","0101","0110","0101","0100","0100","0100","0100","0101","0110","0101","0100","0100","0100","0100","0100","0100","0110","0110","0110","0101","0110","0110","0110","0110","0101","0100","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0101","0101","0101","0110","0101","0011","0101","0101","0011","0100","0101","0100","0011","0011","0010","0010","0010"),
("0011","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0010","0010","0100","0010","0001","0010","0100","0010","0001","0010","0011","0001","0011","0100","0101","0101","0100","0100","0101","0101","1000","1000","0110","0101","0101","0110","0101","0110","0101","0101","0110","0101","0100","0101","0101","0100","0101","0100","0101","0101","0101","0100","0100","0110","0111","0111","0111","0111","0111","0111","0111","0101","0010","0101","0010","0001","0011","0101","0101","0011","0001","0101","0011","0011","0110","0111","0111","0111","0111","0110","0101","0100","0011","0011","0100","0101","0100","0100","0101","0110","0110","0110","0110","0110","0101","0110","0110","0101","0110","0101","0110","0111","0111","0110","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0110","0110","0110","0110","0111","0110","0101","0100","0100","0100","0101","0110","0110","0110","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","1001","1010","1010","1001","1010","1010","0111","0011","0011","0011","0101","0110","0111","0111","0111","1000","0111","0101","0111","0111","0110","0101","0100","0100","0100","0100","0100","0100","0100","0011","0101","0100","0100","0100","0101","0101","0110","0110","0110","0101","0101","0101","0101","0100","0101","0101","0110","0111","0101","0100","0100","0101","0110","0110","0110","0111","0110","0100","0011","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0111","1001","1001","0110","0100","0100","0101","0111","0111","0110","0110","0110","0101","0101","0101","0101","0101","0101","0110","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0011","0101","0111","0101","0100","0100","0110","0101","0101","0100","0100","0011","0011","0101","1000","0110","0110","0110","0110","0111","0111","0110","0110","0111","0111","1000","0100","0010","0001","0001","0101","0100","0011","0010","0001","0011","0100","0011","0100","0011","0011","0011","0001","0010","0011","0010","0010","0011","0011","0011","0100","0011","0010","0001","0000","0011","0011","0100","0101","0001","0010","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0101","0100","0100","0100","0101","0110","0101","0101","0101","0100","0100","0100","0011","0100","0011","0011","0011","0011","0011","0100","0100","0110","1000","0100","0011","0011","0011","0011","0011","0100","0011","0101","0101","0101","0100","0100","0100","0011","0110","1000","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0011","0100","0101","0100","0100","0011","0011","0100","0101","0101","0100","0110","0010","0110","1001","1001","1010","1010","1001","1010","1000","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0101","0101","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0100","0110","0110","0100","0010","0011","0010","0010","0011","0100","0011","0011","0011","0100","0011","0011","0101","0101","0101","0110","0110","0101","0111","1000","1000","0110","0010","0100","1000","0111","0100","0100","0011","0100","0100","0101","0100","0100","0111","1000","0101","0010","0110","1000","0011","0010","0010","0100","0100","0011","0011","0111","0111","0110","0101","0100","0101","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0101","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0010","0010","0010","0001","0010","0010","0100","0011","0011","0010","0010","0100","0101","0011","0100","0101","0101","0101","0100","0100","0101","0101","0100","0100","0100","0011","0011","0110","0110","0110","0110","0101","0110","0110","0110","0110","0101","0101","0110","0111","0110","0110","0111","0110","0110","0110","0110","0110","0101","0101","0110","0110","0101","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010"),
("0011","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0010","0010","0100","0010","0001","0010","0011","0010","0001","0010","0011","0001","0011","0100","0100","0101","0100","0100","0100","0100","0111","1000","0110","0101","0100","0110","0011","0101","0101","0010","0110","0110","0010","0101","0101","0010","0101","0011","0101","0100","0100","0011","0011","0101","0110","0110","0110","0111","0111","0111","0111","0101","0010","0101","0011","0001","0011","0101","0101","0011","0001","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0101","0101","0111","0111","0110","0110","0111","0110","0110","0111","0111","0110","0111","0111","0111","0111","0111","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0110","0110","0101","0101","0101","0101","0110","0011","0101","0101","0011","0101","1000","0111","0110","0110","0110","1000","1000","0111","0111","1001","1010","1010","1000","1000","1010","0111","0100","0100","0100","0101","0110","0111","0111","0111","0111","0111","0101","0101","0110","0101","0101","0100","0100","0100","0101","0110","0110","0011","0011","0100","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0110","0101","0011","0011","0011","0101","0101","0110","0110","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0111","1001","1000","0100","0011","0011","0101","0110","0101","0100","0100","0100","0100","0011","0011","0011","0011","0100","0101","0100","0100","0100","0110","0110","0110","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0101","0100","0011","0011","0100","1000","1000","1000","0111","0111","1000","1000","0110","0101","0101","0100","0110","0101","0101","0011","0010","0101","0100","0011","0010","0001","0010","0011","0011","0101","0100","0101","0100","0011","0011","0100","0011","0011","0101","0100","0100","0101","0011","0001","0001","0000","0011","0011","0101","0101","0010","0011","0100","0100","0100","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0100","0100","0100","0100","0011","0100","0011","0100","0100","0110","0101","0100","0100","0100","0100","0100","0101","0110","0111","0110","0100","0011","0100","0100","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0011","0011","0100","0100","0100","0101","0100","0100","0100","0100","0011","0100","0100","0101","0011","0010","0010","0100","0111","1001","1010","1000","0110","0101","0011","0011","0100","0100","0011","0010","0011","0100","0100","0100","0100","0101","0110","0110","0110","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0110","0101","0100","0100","0100","0101","0100","0101","0100","0101","0101","0101","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0111","0110","0100","0100","0100","0101","0101","0101","0101","0100","0100","0101","0101","0100","0101","0110","0101","0110","0111","0111","1000","1000","1000","1000","0111","0110","0110","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","0011","0010","0010","0100","0111","0111","1000","1000","0110","0101","0100","0011","0100","0100","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0011","0011","0011","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0011","0011","0100","0101","0101","0100","0100","0101","0101","0101","0100","0010","0010","0010","0001","0010","0010","0100","0101","0011","0010","0010","0010","0100","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0011","0100","0111","0110","0110","0110","0101","0110","0110","0101","0110","0100","0100","0110","0111","0101","0101","0110","0110","0101","0100","0101","0110","0101","0011","0011","0100","0100","0011","0011","0010","0011","0011","0010","0010","0011","0010","0011","0011","0010"),
("0011","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0100","0010","0001","0010","0010","0001","0001","0010","0001","0001","0001","0001","0010","0010","0011","0011","0100","0011","0011","0010","0010","0011","0011","0101","0100","0011","0101","0101","0100","0011","0100","0101","0101","0100","0100","0101","0100","0100","0011","0100","0101","0011","0010","0010","0010","0010","0010","0011","0101","0101","0100","0100","0100","0001","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0010","0100","0100","0100","0100","0111","0101","0101","0110","0110","0101","0101","0101","1001","1001","1000","1001","1000","1001","1001","1001","1001","0111","0101","0101","0110","0110","0110","0111","0110","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0110","0101","0101","0110","0111","0111","0110","0110","0110","0111","0110","0101","0101","0110","0110","0111","0111","0111","0110","0110","0111","0011","0101","0110","0011","0010","0110","0111","0101","0101","0100","1000","1000","0101","0110","1001","1010","1000","0100","0100","1001","0111","0011","0011","0011","0100","0101","0101","0101","0110","0111","0111","0111","0110","0100","0100","0100","0100","0100","0011","0011","0101","0110","0011","0010","0011","0101","0101","0110","0110","0110","0110","0110","0100","0010","0101","0110","0110","0110","0101","0101","0111","0110","0110","0110","0110","0111","1000","0111","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0110","1000","0101","0010","0010","0010","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0101","0111","0111","0110","0100","0011","0011","0100","0100","0101","0101","0101","0101","0110","0111","0111","0101","0101","0100","0011","0011","0100","0100","0100","0011","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0101","0101","0101","0101","0101","0100","0100","0101","0100","0100","0100","0100","0101","0101","0100","0011","0110","0100","0011","0011","0001","0011","0100","0011","0110","0101","0110","0101","0100","0100","0100","0011","0100","0101","0100","0100","0101","0011","0001","0001","0000","0011","0011","0101","0101","0011","0011","0100","0100","0011","0011","0011","0100","0101","1000","1000","0111","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0101","0101","0100","0110","0111","1000","0111","1000","0101","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0011","0011","0100","0110","0110","0100","0011","0011","0100","0100","0100","0100","0011","0010","0010","0011","0100","0110","0100","0100","0011","0100","0100","0011","0010","0010","0100","0100","0100","0100","0100","0100","0100","0100","0101","0111","0111","1000","0111","0101","0100","0100","0100","0100","0101","0100","0101","0100","0100","0100","0110","0110","0110","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0100","0101","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0100","0011","0011","0100","0111","0111","1000","1000","0101","0011","0101","0101","0100","0100","0011","0011","0011","0011","0010","0010","0010","0011","0101","0100","0110","0100","0100","0011","0010","0010","0010","0011","0100","0101","0101","0101","0100","0011","0100","0100","0100","0011","0011","0101","1000","1000","0111","0110","0111","0111","0101","0100","0010","0010","0010","0010","0010","0011","0101","0101","0011","0010","0001","0010","0101","0111","0111","0110","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","0101","0110","0110","0101","0110","0110","0110","0110","0100","0100","0110","0111","0110","0110","0110","0101","0100","0011","0100","0101","0101","0011","0011","0100","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010"),
("0100","0011","0011","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0101","0100","0011","0101","0101","0101","0100","0100","0101","0101","0101","0100","0101","0101","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0100","0111","1000","1000","0111","0111","0011","0011","0101","0101","1000","0111","0100","1000","1000","0100","0100","0100","0111","1010","1001","1000","0101","0100","0101","0110","0111","0111","0111","0100","0010","0011","0100","0011","0101","0111","0111","0111","0111","0110","0111","0111","0110","0110","0111","0111","0111","0110","0011","0110","0111","0110","0011","0011","0100","0101","0111","0111","0111","0110","0110","0101","0101","0101","0101","0011","0011","0100","0100","0100","0101","0100","0101","0110","0101","0110","1001","1000","0100","0010","0010","0111","0111","0100","0100","0100","0101","0111","0111","1000","1000","1000","0111","0110","0110","0101","0100","0100","0100","0100","0010","0010","0011","0101","0011","0010","0011","0101","0100","0101","0101","0110","0111","0101","0100","0100","0101","0110","0110","0110","0101","0101","0110","0101","0100","0011","0100","0101","0110","0101","0101","0011","0011","0011","0011","0010","0011","0011","0011","0011","0100","0011","0100","0100","0100","0101","0100","0011","0010","0010","0010","0011","0011","0011","0100","0100","0101","0100","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0011","0100","0100","0100","0101","0100","0101","0100","0101","0111","1000","0110","0101","0100","0010","0010","0100","0101","0100","0011","0100","0100","0100","0101","0100","0100","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0100","0101","0100","0011","0100","0100","0101","0101","0011","0011","0110","0101","0011","0011","0001","0010","0010","0011","0110","0101","0101","0101","0100","0100","0100","0011","0100","0101","0100","0100","0101","0011","0000","0001","0001","0011","0011","0100","0101","0011","0011","0101","0100","0011","0011","0011","0101","0110","0111","0111","0101","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0100","0100","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0101","0101","0101","0110","0110","0110","0110","0101","0101","0101","0111","0111","0101","0110","0110","0101","0101","0100","0110","0111","1000","0101","0110","0110","0101","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0110","0110","0111","0110","0101","0101","0100","0100","0100","0101","0101","0100","0100","0011","0100","0100","0011","0011","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0010","0010","0100","0100","0100","0100","0101","0101","0100","0100","0100","0101","0110","0110","0101","0100","0011","0100","0011","0100","0100","0011","0011","0011","0011","0011","0110","0110","0110","0111","1000","0101","0101","1000","0111","0100","0110","1000","0110","0101","0111","1000","0111","0110","0110","0110","0110","0110","0101","0101","0010","0010","0101","1000","1000","1000","0111","0100","0101","1000","0111","0110","0101","0101","0101","0101","0101","0101","0101","0111","1000","0101","0011","0110","1000","0011","0010","0010","0011","0100","0011","0011","0110","0110","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0100","0110","0101","0111","0111","0111","0101","0010","0010","0010","0011","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0011","0100","0110","0111","0111","0110","0111","0111","0110","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0001","0010","0101","0111","0111","0101","0011","0011","0011","0011","0011","0011","0011","0100","0010","0010","0011","0111","0110","0110","0110","0101","0110","0110","0110","0101","0101","0100","0101","0110","0110","0101","0100","0100","0101","0101","0100","0101","0101","0011","0011","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010"),
("0100","0011","0011","0010","0010","0010","0010","0011","0100","0100","0100","0100","0101","0100","0100","0100","0011","0100","0101","0110","0101","0110","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0110","0101","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0110","0101","0101","0101","0101","0110","0110","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0110","0110","0110","0110","0101","0100","0100","0100","0101","0110","0110","0101","0101","0101","0100","0101","0110","0111","1001","1001","0111","0100","0011","0011","0100","0101","0110","0110","0011","0010","0010","0011","0011","0101","0111","0111","0111","0101","0100","0100","0100","0101","0101","0101","0101","0101","0100","0011","0101","0110","0110","0100","0101","0101","0101","0110","0110","0110","0110","0101","0101","0110","0101","0101","0110","0101","0101","0101","0101","0101","0110","0111","0111","0101","0101","0110","0100","0010","0010","0010","0100","0111","0011","0011","0011","0100","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0010","0010","0010","0010","0011","0010","0010","0010","0100","0100","0100","0101","0110","0110","0100","0100","0110","0110","0110","0101","0110","0101","0100","0101","0100","0011","0011","0011","0100","0011","0011","0011","0010","0011","0010","0010","0011","0011","0100","0100","0100","0100","0101","0101","0110","0110","0101","0101","0011","0010","0011","0011","0011","0011","0011","0100","0101","0101","0100","0100","0100","0100","0100","0101","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0010","0010","0011","0110","0111","0110","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","0111","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0110","0110","0101","0011","0011","0110","0101","0011","0011","0001","0001","0001","0011","0110","0101","0101","0100","0011","0100","0100","0011","0100","0101","0100","0100","0101","0011","0001","0001","0001","0011","0011","0100","0101","0011","0011","0100","0100","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0011","0010","0010","0011","0100","0100","0100","0100","0100","0101","0110","0101","0111","0110","0110","0110","0101","0101","0101","0111","0110","0111","1000","1000","0111","0110","0101","0110","0111","1000","0110","0111","0110","0101","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0110","0110","0111","0110","0110","0101","0001","0010","0011","0110","0100","0010","0010","0001","0100","0100","0010","0011","0010","0010","0011","0011","0100","0101","0110","0110","0110","0110","0100","0010","0010","0011","0101","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0011","0100","0100","0100","0011","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0110","0110","0111","0111","0011","0011","1000","0110","0001","0100","0110","0100","0010","0111","1000","0100","0010","0010","0100","0011","0011","0010","0010","0010","0010","0010","0111","1000","1000","0110","0011","0100","1000","0111","0101","0101","0101","0100","0100","0100","0100","0100","0111","1000","0101","0011","0110","1000","0011","0010","0010","0011","0100","0100","0100","0111","0101","0100","0101","0100","0100","0101","0110","0110","0111","0101","0101","0110","0101","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0100","0100","0110","0110","0111","1000","0111","0011","0010","0010","0010","0010","0010","0010","0010","0100","0100","0010","0010","0010","0011","0100","0100","0100","0011","0100","0011","0011","0011","0011","0011","0100","0010","0010","0011","0111","0110","0110","0110","0101","0110","0101","0100","0100","0011","0011","0100","0100","0101","0100","0100","0100","0100","0101","0101","0101","0101","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0100","0100","0011","0010","0010","0010","0010","0011","0011","0100","0011","0100","0011","0011","0011","0011","0011","0100","0110","0101","0011","0100","0110","0101","0011","0011","0101","0101","0100","0100","0101","0101","0110","0110","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0110","0110","0111","1000","0110","0101","0110","0110","0110","0101","0111","0111","0101","0100","0100","0011","0010","0010","0011","0100","0100","0110","0111","0100","0110","1000","0111","0101","0011","0101","1000","0111","0100","0110","0111","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0100","0100","1000","1000","1001","1000","1001","1001","1001","0111","0100","0011","0011","0100","0100","0011","0010","0010","0010","0010","0011","0100","0110","0110","0110","0101","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0111","0111","0111","0111","0110","0110","0110","0110","0110","0101","0110","0111","0110","0101","0111","0110","0101","0110","0110","0110","0110","0110","0110","0101","0101","0011","0010","0010","0010","0010","0011","0110","0100","0011","0011","0100","0101","0101","0100","0101","0101","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0110","0101","0111","0110","0011","0011","0101","0110","0110","0101","0111","0110","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0101","0101","0101","0110","0101","0101","0110","0110","0110","0110","0111","0101","0101","0100","0100","0100","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0011","0011","0100","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0100","0011","0100","0100","0101","0101","0101","0010","0010","0010","0011","0101","0101","0101","0110","0111","0111","0110","0101","0111","0111","0111","0111","0111","1000","0101","0101","0110","0100","0101","0110","0111","0100","0101","0110","0100","0101","0110","0101","0100","0101","0101","0011","0011","0110","0101","0011","0011","0001","0011","0100","0100","0101","0101","0101","0100","0011","0100","0100","0011","0100","0101","0100","0100","0101","0011","0010","0010","0001","0011","0011","0100","0101","0011","0011","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0010","0010","0011","0100","0101","0101","0101","0100","0101","0110","0101","0111","0111","0111","0110","0111","0111","0110","0101","0101","0101","0111","0110","0101","0101","0100","0110","0111","0110","0101","0100","0100","0101","0110","0101","0100","0110","0111","1000","0111","0101","0100","0100","0100","0100","0100","0101","0101","0110","0101","0101","0101","0010","0010","0011","0110","0100","0010","0010","0010","0100","0100","0011","0100","0011","0010","0011","0100","0100","0101","0110","0110","0101","0100","0100","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0010","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0110","0110","0110","0110","0110","0100","0100","0111","0101","0100","0101","0110","0101","0100","0110","0110","0111","0111","0111","0111","0111","0111","0111","0011","0010","0010","0011","0111","0111","1000","0111","0110","0111","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","0111","0111","1000","0100","0010","0010","0100","0111","1000","1000","1000","0110","0100","0101","0110","0110","0110","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","1000","0111","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0010","0010","0010","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0100","0101","0110","0101","0101","0100","0100","0100","0011","0011","0011","0011","0010","0011","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0110","0101","0011","0010","0010","0010","0010","0011","0011","0011","0100","0100","0011","0011","0011","0010","0010","0011","0110","0011","0010","0010","0100","0100","0010","0011","0101","0100","0100","0100","0011","0011","0100","0100","0011","0100","0011","0011","0100","0101","0101","0101","0101","0110","0111","0110","0111","1000","0111","0110","0110","0111","0111","0110","0111","0111","0100","0100","0011","0011","0010","0010","0011","0011","0011","0110","0101","0011","0100","0111","0110","0011","0010","0011","0111","0110","0010","0100","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","0011","0011","0110","1000","1000","0111","1000","1001","1001","1000","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0101","0100","0011","0011","0011","0011","0101","0110","0101","0011","0011","0100","0011","0011","0101","0110","0110","0100","0101","0101","0101","0100","0010","0010","0010","0010","0011","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0100","0100","0010","0010","0100","0101","0110","0101","0110","0110","0101","0101","0100","0011","0010","0011","0101","0110","0101","0100","0110","0110","0110","0111","0110","0110","0110","0111","1000","0111","0101","0011","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0101","0110","0110","0110","0110","0101","0101","0101","0100","0100","0100","0100","0100","0101","0100","0011","0100","0100","0101","0110","0101","0010","0010","0010","0010","0010","0011","0100","0110","0100","0101","0111","0101","0110","0110","0101","0110","0110","1000","0110","0110","0101","0011","0011","0100","0110","0101","0101","0110","0110","0110","0110","0110","0101","0101","0101","0011","0011","0110","0101","0011","0011","0010","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0011","0100","0101","0101","0100","0101","0011","0010","0010","0001","0011","0011","0100","0110","0011","0011","0101","0100","0101","0100","0101","0101","0100","0100","0100","0100","0100","0100","0011","0100","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0100","0011","0011","0010","0010","0011","0101","0101","0101","0100","0101","0110","0101","0111","0111","0101","0101","0110","0111","0110","0111","0110","0101","0100","0100","0101","0101","0100","0101","0110","0101","0011","0100","0101","0101","0110","0101","0101","0101","0110","0111","0111","0101","0100","0100","0011","0100","0100","0101","0101","0101","0101","0101","0101","0011","0011","0011","0101","0100","0011","0100","0011","0100","0100","0011","0110","0110","0100","0100","0100","0100","0101","0101","0110","0101","0100","0100","0101","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0011","0100","0100","0100","0100","0101","0101","0100","0011","0011","0011","0100","0100","0100","0010","0011","0100","0011","0011","0011","0011","0011","0100","0110","0110","0110","0110","0110","0110","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","0100","0011","0010","0010","0011","0100","0110","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","0111","1000","1000","0100","0011","0011","0100","0111","0111","0111","1000","0101","0011","0101","0101","0101","0110","0111","0111","0110","0111","1000","1000","1000","0111","0110","0110","0110","0111","1000","1000","1000","1000","1000","0111","0110","0110","0011","0011","0011","0100","0100","0100","0011","0011","0100","0011","0011","0011","0011","0100","0101","0110","0100","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0100","0100","0101","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0100","0100","0011","0010","0010","0010","0010","0010","0011","0011","0100","0100","0011","0011","0011","0010","0010","0011","0110","0011","0010","0010","0100","0100","0010","0011","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0101","0100","0100","0011","0011","0100","0100","0101","0110","0101","0011","0011","0111","0111","0011","0010","0011","0111","0101","0001","0100","0110","0110","0111","1000","0111","0111","1000","1000","1000","1000","0111","0110","0011","0011","0011","0110","0111","0101","0111","1000","1000","0111","0100","0100","0101","0100","0100","0011","0010","0010","0010","0011","0100","0101","0100","0011","0100","0100","0011","0010","0100","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0100","0010","0010","0010","0011","0100","0101","0101","0011","0011","0100","0011","0011","0101","0110","0110","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0011","0101","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0011","0010","0010","0011","0101","0101","0110","0101","0110","0111","0110","0100","0011","0010","0010","0100","0101","0011","0011","0011","0011","0100","0100","0011","0100","0110","0111","1000","0110","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0110","0101","0110","0111","0110","0101","0101","0101","0101","0100","0011","0100","0100","0011","0011","0011","0100","0100","0101","0100","0011","0010","0010","0010","0010","0101","0110","0110","0100","0110","1000","1000","1000","1001","1001","1001","1001","1001","0111","0110","0100","0010","0010","0011","0011","0100","0101","0101","0100","0011","0101","0111","0111","0110","0101","0011","0011","0101","0101","0011","0010","0010","0011","0100","0100","0101","0101","0101","0100","0100","0100","0100","0011","0100","0101","0101","0100","0101","0011","0010","0010","0001","0011","0011","0100","0110","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0110","0101","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0100","0101","0100","0011","0011","0010","0010","0011","0100","0101","0101","0101","0101","0101","0110","0111","0100","0101","0101","0100","0101","0101","0101","0111","0110","0100","0011","0011","0011","0101","0101","0100","0100","0100","0100","0101","0100","0100","0101","0101","0101","0100","0101","0110","0110","0110","0101","0101","0100","0100","0101","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0101","0100","0101","0101","0100","0010","0100","0100","0100","0100","0101","0101","0101","0110","0110","0110","0101","0100","0101","0100","0010","0010","0011","0100","0100","0100","0011","0100","0100","0011","0010","0010","0010","0010","0100","0100","0100","0100","0100","0011","0011","0011","0010","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0110","0110","0110","0110","0111","0111","0101","0110","0111","0101","0111","1000","0111","0110","0110","0110","1000","0101","0011","0111","1000","0101","0010","0010","0010","0010","0010","0100","0110","0111","0110","0011","0101","1000","0111","0101","0101","0100","0101","0101","0100","0100","0100","0111","1000","0101","0011","0110","1000","0100","0011","0011","0100","0100","0011","0011","0110","0101","0010","0101","0101","0100","0110","0111","0111","0100","0101","1000","0111","1000","0111","0101","0100","0101","1000","0111","1000","1000","1000","1000","0101","0011","0011","0011","0011","0011","0100","0101","0101","0101","0101","0101","0100","0010","0011","0011","0011","0011","0101","0101","0100","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0011","0100","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0011","0011","0100","0010","0010","0010","0010","0010","0011","0100","0100","0011","0011","0010","0011","0010","0010","0011","0110","0011","0010","0010","0100","0101","0010","0011","0011","0011","0011","0100","0100","0100","0011","0010","0011","0011","0011","0010","0010","0011","0101","0101","0101","0111","0111","0110","0110","0110","0110","0110","0110","0111","1000","1000","1000","0110","0101","0101","0100","0100","0100","0100","0011","0100","0101","0110","0101","0010","0011","0111","0110","0011","0011","0011","0111","0101","0001","0011","0110","0111","1000","1000","1000","1000","1000","1000","0111","1000","0110","0011","0011","0010","0011","0101","0111","0101","0111","1000","1000","0110","0110","0110","0101","0100","0101","0011","0010","0010","0010","0011","0100","0101","0101","0100","0100","0100","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0100","0101","0101","0011","0101","0101","0101","0101","0110","0110","0111","0110","0101","0101","0100","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0011","0101","0101","0100","0100","0100","0100","0100","0100","0101","0100","0100","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0100","0100","0011","0010","0011","0100","0101","0100","0100","0110","0101","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0101","0110","0110","0101","0101","0110","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0110","1000","0101","0101","0101","0101","0110","0100","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0110","0110","0110","0100","0101","0110","0101","0110","0110","0110","0110","0110","1000","0110","0100","0011","0100","0011","0011","0011","0100","0110","0110","0011","0100","0101","0110","0110","0110","0110","0100","0011","0101","0100","0011","0011","0010","0011","0011","0011","0101","0101","0110","0101","0100","0100","0100","0011","0100","0101","0101","0101","0101","0011","0001","0001","0001","0011","0011","0101","0110","0011","0011","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0011","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0011","0011","0100","0100","0101","0101","0100","0011","0011","0010","0010","0010","0011","0100","0101","0101","0101","0101","0100","0101","0011","0011","0101","0101","0101","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0101","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0100","0010","0010","0010","0011","0101","0010","0011","0100","0011","0010","0011","0100","0011","0011","0100","0100","0100","0101","0101","0101","0100","0011","0100","0100","0010","0010","0011","0100","0100","0100","0011","0100","0011","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0010","0010","0010","0010","0011","0011","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0110","0110","0110","0110","0110","0100","0100","0100","0100","0101","0101","0100","0010","0010","0011","0111","0101","0011","0111","0111","0100","0010","0010","0010","0010","0010","0011","0100","0111","0110","0011","0101","1000","0111","0100","0100","0100","0100","0101","0100","0100","0100","0111","1000","0101","0011","0110","1000","0100","0011","0011","0100","0101","0101","0101","0111","0100","0001","0100","0101","0100","0110","0111","1000","0101","0101","1000","0111","1000","0110","0101","1000","0111","0111","1000","1000","1000","1000","1000","0111","0111","0110","0100","0011","0011","0100","0100","0100","0100","0101","0101","0100","0011","0011","0100","0100","0101","0101","0011","0010","0010","0010","0010","0010","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0011","0011","0011","0010","0010","0010","0010","0011","0100","0011","0011","0011","0010","0010","0011","0011","0010","0011","0110","0011","0010","0011","0100","0101","0010","0011","0011","0100","0011","0010","0011","0101","0101","0011","0100","0011","0011","0011","0011","0100","0110","0110","0101","0110","0111","0111","1000","1000","1000","0111","0111","0110","0111","0111","1000","0110","0101","0101","0100","0100","0100","0101","0100","0100","0100","0110","0101","0011","0100","0111","0111","0100","0100","0011","0111","0110","0011","0100","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","0110","0011","0010","0010","0011","0011","0100","0100","0110","1000","1000","0100","0101","0101","0101","0101","0011","0010","0010","0010","0010","0011","0011","0100","0110","0101","0101","0100","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0101","0110","0110","0110","0110","0110","0100","0011","0011","0011","0011","0100","0100","0100","0011","0100","0110","0110","0111","1000","1000","1000","1000","0111","0111","0101","0011","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0101","0110","0101","0101","0100","0100","0110","0101","0101","0110","0101","0110","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0110","0100","0010","0011","0100","0101","0100","0101","0111","0101","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0101","0100","0101","0101","0110","0101","0101","0101","0100","0101","0101","0011","0011","0100","0101","0100","0101","0110","0110","0101","0101","0101","0101","0101","0101","0110","0111","0101","0100","0110","0101","0101","0101","0100","0110","0100","0100","0100","0100","0110","0111","0110","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0110","0101","0100","0100","0111","0110","0110","0101","0101","0110","0110","1000","0111","0100","0100","0011","0011","0011","0011","0100","0101","0101","0100","0100","0101","0111","0101","0101","0101","0100","0100","0110","0101","0011","0011","0010","0100","0100","0011","0110","0101","0101","0100","0100","0100","0100","0011","0011","0100","0100","0101","0101","0011","0010","0010","0001","0011","0011","0100","0110","0101","0011","0100","0101","1000","0111","0101","0101","0101","0100","0101","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0011","0010","0010","0010","0010","0100","0100","0100","0101","0100","0100","0011","0010","0010","0100","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0100","0010","0010","0010","0011","0101","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0100","0100","0011","0010","0010","0010","0010","0011","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0100","0100","0011","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0011","0011","0010","0010","0011","0011","0011","0100","0101","0110","0110","0101","0101","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0011","0110","0100","0100","0101","0101","0011","0010","0010","0010","0010","0010","0010","0011","0111","0111","0110","0111","1000","1000","1000","1000","1000","1000","0110","0111","0110","0111","0111","0111","0111","0111","1000","1000","0100","0011","0100","0100","0111","1000","1000","0111","0011","0010","0011","0011","0100","0110","0111","1000","0101","0101","0111","0111","0111","0101","0011","0110","0111","0111","1000","0111","0111","0110","0111","0111","0110","0101","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0101","0011","0010","0010","0010","0010","0010","0011","0100","0100","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0110","0011","0010","0010","0011","0100","0010","0011","0011","0010","0010","0011","0101","0110","0101","0011","0100","0101","0100","0011","0010","0011","0100","0100","0100","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0101","0100","0101","0101","0101","0101","0101","0101","0100","0110","0101","0011","0011","0111","0111","0100","0011","0011","0110","0110","0011","0100","0111","1000","0111","1000","0111","1000","0111","1000","1000","0101","0100","0011","0010","0010","0010","0011","0011","0011","0110","1000","0111","0011","0100","0101","0110","0101","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0100","0100","0100","0010","0011","0110","1000","1000","1001","1000","1000","1000","0111","1000","0101","0011","0010","0010","0010","0011","0100","0100","0100","0100","0101","0101","0011","0011","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0110","0101","0100","0011","0101","0101","0101","0110","0110","0110","0101","0100","0011","0010","0011","0111","0100","0101","0101","0100","0011","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0011","0011","0100","0100","0100","0101","0110","0110","0101","0110","0101","0110","0110","0110","0110","0101","0110","0101","0110","0101","0110","0101","0110","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0111","0110","0110","0110","0101","0100","0100","0100","0101","0100","0101","0111","0110","0101","0110","0111","0110","0111","0110","0011","0100","0011","0011","0010","0011","0100","0100","0101","0100","0011","0101","0101","0011","0100","0101","0100","0110","0110","0100","0011","0011","0010","0011","0011","0011","0110","0101","0100","0100","0011","0011","0100","0011","0011","0100","0100","0101","0101","0011","0010","0010","0001","0011","0011","0100","0110","0101","0011","0100","0101","0111","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0011","0010","0010","0010","0010","0010","0011","0011","0011","0101","0100","0100","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0100","0011","0010","0010","0010","0010","0010","0011","0100","0011","0011","0011","0100","0101","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0010","0010","0011","0010","0010","0011","0100","0100","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0100","0101","0100","0101","0100","0100","0100","0100","0011","0100","0100","0100","0100","0011","0011","0011","0100","0011","0100","0100","0011","0010","0010","0010","0010","0010","0011","0100","0100","0101","0100","0101","0101","0101","1000","1000","1000","0101","0101","0101","0101","0101","0110","0110","0111","0111","1000","0100","0011","0100","0100","0110","0111","0110","0100","0011","0001","0010","0011","0100","0110","0111","0111","0101","0101","0110","0110","0110","0011","0010","0100","0110","0111","0111","0101","0110","0100","0101","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0100","0100","0011","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0110","0011","0010","0010","0011","0100","0010","0011","0100","0011","0011","0100","0101","0101","0101","0100","0100","0100","0100","0011","0010","0011","0100","0100","0101","0111","1000","1000","0111","0101","0111","1000","1000","1000","1000","0111","0111","0110","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0010","0011","0111","0111","0011","0010","0010","0110","0110","0010","0011","0111","1000","1000","0111","1000","0111","1000","1000","1000","0111","0101","0011","0010","0010","0011","0100","0011","0100","0110","1000","0111","0100","0011","0100","0100","0101","0100","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0100","0011","0011","0011","0010","0101","0110","1000","1001","1001","1001","1000","0111","1000","0111","0011","0010","0010","0010","0100","0100","0100","0100","0100","0101","0100","0011","0010","0100","0101","0101","0100","0101","0101","0110","0110","0110","0101","0110","0101","0100","0100","0101","0100","0101","0110","0110","0101","0101","0101","0101","0110","0111","0100","0010","0010","0011","0101","0100","0100","0011","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0101","0101","0100","0100","0100","0101","0101","0101","0100","0100","0010","0100","0110","0110","0110","0011","0101","0011","0100","0100","0011","0101","0011","0101","0010","0101","0010","0101","0011","0100","0100","0100","0111","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0011","0100","0101","0011","0010","0010","0011","0010","0010","0011","0011","0100","0101","0100","0011","0101","0100","0010","0100","0100","0100","0101","0110","0101","0011","0011","0001","0010","0001","0011","0110","0101","0101","0100","0011","0100","0100","0011","0011","0100","0100","0101","0101","0011","0001","0001","0001","0011","0011","0101","0110","0101","0011","0101","0100","0100","0011","0100","0100","0100","0011","0011","0011","0100","0100","0100","0011","0110","0101","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0011","0100","0100","0011","0010","0010","0010","0011","0100","0100","0100","0011","0011","0100","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0101","0101","0101","0101","0100","0101","0100","0101","0100","0100","0100","0100","0011","0100","0011","0011","0011","0011","0011","0100","0011","0100","0100","0100","0100","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0011","0011","0100","0011","0011","0011","0100","0100","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0100","0100","0011","0011","0011","0011","0100","0101","0101","0101","0101","0101","0101","0110","0101","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0011","0011","0011","0011","0100","0101","0100","0010","0101","1000","0100","0011","0100","0100","0100","0100","0011","0010","0010","0010","0010","0011","0011","0101","0111","0111","0100","0100","0101","0101","0101","0011","0010","0011","0100","0110","0101","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0101","0100","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0010","0010","0011","0110","0011","0010","0010","0011","0100","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0111","0111","1000","0100","0001","0011","0111","1000","1000","1000","1000","0111","0110","0100","0101","0101","0101","0101","0101","0101","0110","0101","0110","0101","0011","0011","0111","0111","0011","0011","0011","0111","0110","0010","0011","0111","1000","1000","1000","1000","1000","1000","1000","0111","0101","0100","0011","0010","0010","0011","0100","0100","0100","0110","1000","1000","0100","0100","0100","0101","0101","0100","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0100","0011","0011","0011","0100","0101","0110","0110","0110","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0101","0110","0111","1000","1000","1000","0111","1000","0101","0010","0010","0010","0010","0100","0101","0101","0101","0100","0101","0011","0010","0010","0011","0101","0101","0100","0101","0110","0110","0110","0111","0110","0110","0110","0100","0100","0101","0100","0101","0111","0111","0101","0101","0101","0011","0101","0111","0100","0010","0010","0010","0100","0100","0100","0011","0010","0010","0101","0110","0110","0101","0110","0110","0110","0101","0101","0101","0110","0110","0101","0101","0100","0010","0100","0100","0100","0101","0100","0101","0100","0010","0100","0101","0110","0111","0011","0101","0100","0101","0100","0100","0101","0011","0101","0010","0101","0011","0101","0011","0100","0100","0100","0111","0100","0010","0011","0011","0011","0011","0010","0010","0011","0010","0010","0011","0100","0101","0100","0110","0111","0101","0011","0011","0100","0011","0100","0100","0011","0011","0100","0100","0011","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0101","0101","0100","0110","0111","0101","0011","0011","0001","0010","0010","0011","0110","0110","0110","0101","0100","0100","0101","0100","0100","0101","0101","0101","0110","0011","0001","0001","0001","0011","0100","0101","0110","0110","0100","0101","0100","0100","0011","0011","0100","0100","0011","0011","0011","0100","0100","0100","0011","0101","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0100","0011","0100","0100","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0101","0101","0110","0101","0100","0101","0100","0101","0100","0100","0100","0100","0011","0011","0011","0100","0100","0011","0100","0100","0100","0100","0010","0010","0011","0101","0100","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0100","0100","0011","0101","1000","0100","0011","0100","0100","0110","0110","0110","0100","0010","0010","0010","0010","0011","0101","0111","0111","0100","0011","0100","0100","0100","0011","0010","0010","0100","0101","0101","0100","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0101","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0100","0101","0101","0011","0010","0010","0011","0101","0011","0010","0010","0011","0100","0011","0011","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0011","0011","0100","0101","0111","0111","0111","0011","0001","0010","0111","1000","1000","1000","1000","1000","0110","0100","0110","0110","0110","0101","0101","0110","0110","0110","0110","0101","0011","0011","0111","0110","0011","0011","0011","0111","0110","0001","0011","0111","0111","1000","1000","1000","1000","1000","0111","0110","0100","0011","0010","0010","0010","0010","0010","0010","0011","0110","1000","0111","0100","0011","0100","0011","0011","0100","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0110","0110","0101","0100","0011","0011","0100","0100","0100","0101","0101","0100","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0100","0011","0010","0010","0010","0010","0011","0011","0100","0100","0011","0101","0100","0011","0010","0011","0101","0111","0110","0101","0101","0110","0110","0111","0110","0111","1000","0110","0100","0111","0101","0100","0100","0101","0101","0101","0101","0011","0100","0101","0011","0010","0010","0010","0100","0011","0011","0011","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0010","0010","0011","0011","0100","0100","0100","0100","0010","0100","0101","0111","0111","0011","0101","0100","0101","0100","0100","0101","0011","0110","0011","0101","0011","0101","0100","0100","0101","0100","0111","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0101","0011","0110","0111","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0011","0100","0101","0110","0100","0110","0111","0110","0011","0011","0001","0010","0010","0011","0110","0110","0101","0101","0100","0100","0101","0100","0100","0101","0101","0101","0110","0011","0001","0001","0000","0011","0011","0101","0110","0110","0100","0101","0101","0100","0100","0100","0100","0100","0011","0011","0100","0100","0011","0011","0011","0011","0100","0111","0111","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0101","1000","0011","0011","0011","0011","0011","0011","0011","0011","0110","0110","0100","0100","0101","0011","0010","0100","0100","0101","0101","0011","0011","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0100","0011","0011","0011","0011","0100","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0011","0011","0100","0100","0011","0011","0101","0101","0011","0011","0011","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0100","0100","0100","0101","0111","0100","0100","0100","0100","0110","0111","0101","0011","0010","0010","0010","0010","0011","0100","0110","0101","0100","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0101","0100","0010","0010","0011","0011","0011","0011","0010","0011","0101","0110","0110","0110","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0011","0100","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0100","0101","0101","0110","0110","0111","1000","0011","0010","0011","0111","0111","0110","1000","1000","1000","0110","0101","0110","0110","0101","0100","0100","0100","0100","0101","0110","0111","0110","0110","1000","0111","0110","0110","0110","0111","0111","0110","0111","0101","0100","0110","1000","1000","1000","1000","1000","0110","0011","0010","0010","0010","0010","0010","0010","0010","0011","0110","1000","0111","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0101","0100","0100","0101","0101","0011","0011","0011","0100","0101","0101","0101","0101","0011","0010","0010","0011","0101","0101","0101","0101","0101","0101","0101","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0100","0011","0010","0011","0100","0101","0101","0100","0011","0101","0111","0111","0111","0110","0110","0110","0100","0101","0100","0100","0110","0110","0100","0101","0101","0011","0101","0100","0010","0010","0010","0010","0010","0011","0011","0011","0010","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0100","0110","0111","0100","0101","0100","0110","0101","0100","0101","0011","0110","0011","0101","0100","0101","0100","0100","0101","0100","0111","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0110","0101","0110","0111","0100","0010","0010","0011","0010","0010","0011","0010","0011","0100","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0110","0100","0110","0111","0110","0011","0011","0001","0010","0010","0011","0110","0110","0110","0101","0100","0100","0101","0100","0100","0101","0101","0101","0110","0100","0001","0001","0000","0011","0100","0101","0110","0101","0100","0101","0110","0111","0110","0110","0101","0100","0100","0100","0011","0011","0011","0010","0011","0011","0100","0101","0110","0111","1000","1000","1000","1000","0111","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0110","0110","0101","0011","0010","0011","0011","0110","0101","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0010","0010","0010","0011","0100","0100","0100","0011","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0100","0011","0011","0011","0011","0010","0011","0011","0011","0100","0101","0011","0011","0011","0011","0100","0110","0100","0010","0010","0010","0010","0010","0010","0011","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010"),
("0100","0011","0011","0011","0100","0010","0010","0010","0011","0100","0110","0110","0110","0101","0101","0101","0101","0101","0101","0110","0011","0100","0101","0100","0011","0100","0100","0011","0011","0011","0010","0011","0011","0010","0010","0010","0011","0011","0011","0100","0101","0101","0101","0101","0101","1000","0011","0011","0011","0111","0110","0011","0111","1000","1000","0110","0101","0110","0101","0100","0011","0011","0011","0010","0011","0110","1001","1001","1001","1000","1000","0111","0101","1000","1000","1000","1000","1000","0110","0011","0011","0101","0111","0110","0111","1000","0101","0100","0011","0010","0010","0010","0010","0011","0011","0011","0101","1000","1000","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0101","0101","0101","0101","0100","0011","0010","0010","0011","0100","0101","0101","0101","0100","0100","0100","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0100","0011","0010","0101","0111","0111","0111","0110","0100","0101","0101","0101","0100","0101","0111","0110","0100","0101","0101","0011","0100","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0111","0100","0101","0100","0101","0101","0101","0110","0011","0110","0011","0101","0100","0101","0100","0100","0101","0100","0111","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0110","0111","0111","0111","0100","0010","0010","0010","0011","0010","0011","0011","0010","0011","0100","0010","0001","0010","0010","0010","0001","0010","0010","0010","0011","0100","0100","0100","0011","0100","0100","0011","0011","0011","0101","0110","0100","0101","0110","0101","0011","0011","0001","0010","0010","0011","0101","0110","0110","0101","0100","0100","0100","0011","0100","0100","0101","0101","0101","0011","0001","0010","0001","0011","0100","0100","0101","0100","0100","0101","0101","0110","0101","0101","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0100","0101","0101","0101","0101","0101","0110","0111","0110","0110","0111","0111","1000","1000","1000","1001","1001","1010","1000","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","0111","0100","0010","0010","0010","0010","0100","0100","0010","0011","0100","0100","0100","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0101","0101","0011","0100","0100","0011","0100","0011","0011","0011","0100","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0100","0100","0101","0101","0011","0011","0100","0100","0011","0011","0010","0011","0011","0011","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0101","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0011","0011","0010","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0011","0011","0010","0010","0001","0001","0001","0010","0010"),
("0011","0100","0101","0101","0101","0100","0011","0010","0011","0101","0110","0110","0110","0110","0100","0101","0110","0100","0101","0101","0010","0010","0101","0100","0011","0100","0100","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0100","0100","0011","0100","0100","0101","0101","0101","1000","0011","0011","0011","0111","0110","0011","0111","1000","1000","0110","0101","0101","0100","0011","0011","0011","0010","0010","0010","0101","1000","1000","1001","1000","1000","0111","0010","0111","1000","1000","1000","1001","0110","0010","0011","0100","0100","0101","0111","0101","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0100","0100","0100","0011","0010","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0010","0010","0010","0100","0100","0101","0101","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0100","0011","0010","0100","0111","0111","0111","0111","0011","0100","0111","1000","0101","0100","0011","0100","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0101","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0100","0110","0100","0101","0100","0100","0101","0101","0110","0011","0110","0011","0101","0100","0101","0101","0100","0101","0100","0111","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0101","0101","0110","0111","0101","0100","0100","0101","0101","0101","0101","0101","0100","0101","0101","0011","0010","0010","0011","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0010","0010","0011","0011","0101","0101","0100","0100","0101","0101","0100","0011","0001","0010","0010","0010","0101","0110","0110","0101","0100","0100","0011","0011","0011","0100","0100","0101","0100","0011","0001","0001","0000","0011","0100","0100","0100","0100","0011","0101","0100","0100","0100","0011","0010","0100","0011","0100","0100","0100","0100","0011","0011","0100","0100","0101","0101","0110","0110","0110","0101","0101","0100","0100","0100","0110","0110","0101","0100","0100","0101","1000","0111","0100","0100","0100","0100","0100","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0100","0100","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0010","0011","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0100","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0100","0011","0010","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","0100","0011","0010","0010","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0101","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0011","0011","0011","0011","0011","0100","0011","0110","0110","0010","0011","0100","0011","0010","0010","0101","0101","0011","0010","0010","0010","0011","0011","0011","0011","0010","0011","0101","0100","0011","0011","0100","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0001","0001","0010","0010"),
("0101","0101","0101","0110","0110","0110","0011","0010","0011","0100","0011","0010","0010","0010","0100","0101","0101","0101","0101","0110","0010","0011","0101","0100","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0101","0101","0110","0100","0101","1000","0011","0010","0011","0111","0110","0011","0111","1000","1000","0111","0101","0100","0011","0011","0011","0010","0010","0010","0010","0101","1000","1000","1000","1000","1000","0111","0010","0111","1000","1001","1000","1001","0101","0010","0011","0011","0010","0011","0100","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0110","0101","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0011","0100","0100","0100","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0100","0011","0011","0011","0010","0011","0101","0111","0111","0110","0011","0011","0100","0110","0101","0101","0101","0101","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0101","0101","0100","0101","0101","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0111","0100","0101","0101","0101","0101","0100","0110","0011","0110","0011","0101","0100","0101","0101","0100","0110","0100","0111","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0101","0011","0110","0111","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0011","0010","0011","0011","0011","0101","0110","0100","0101","0111","0110","0100","0100","0001","0001","0010","0010","0110","0110","0110","0101","0011","0100","0011","0011","0100","0100","0100","0101","0101","0011","0001","0010","0010","0011","0100","0100","0101","0101","0011","0101","0101","0100","0100","0100","0011","0100","0011","0011","0011","0011","0100","0100","0101","0100","0100","0100","0110","0110","0110","0101","0101","0100","0100","0011","0011","0100","0100","0011","0010","0010","0011","0100","0101","0100","0100","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0101","0100","0011","0011","0011","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0100","0100","0100","0010","0010","0101","0101","0101","0101","0101","0110","0110","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0011","0100","0011","0011","0011","0011","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0100","0100","0011","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0010","0100","0011","0011","0011","0100","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0100","0011","0011","0111","0111","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0101","0100","0100","0100","0100","0011","0010","0011","0011","0011","0011","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0011","0011","0010","0010","0010","0010","0001","0010","0010"),
("0110","0101","0101","0101","0101","0101","0101","0100","0011","0100","0100","0011","0010","0010","0100","0101","0110","0100","0101","0110","0101","0100","0101","0100","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0100","0101","0110","0110","0100","0101","1000","0100","0010","0011","0111","0110","0011","0111","1000","1000","0111","0101","0100","0011","0011","0010","0010","0010","0001","0001","0101","1000","1001","1000","1000","1000","1000","0111","1000","1001","1001","1001","1001","0110","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0100","0100","0110","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0010","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0111","0101","0010","0010","0100","0101","0101","0101","0111","0110","0100","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0100","0100","0101","0101","0100","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0011","0111","0100","0101","0101","0101","0101","0011","0110","0011","0110","0011","0101","0100","0101","0101","0100","0110","0100","0111","0100","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0101","0100","0110","0111","0110","0101","0101","0101","0101","0011","0100","0100","0100","0010","0100","0101","0101","0101","0100","0101","0101","0100","0110","0110","0110","0101","0100","0100","0100","0100","0011","0011","0011","0011","0101","0110","0100","0101","0110","0110","0101","0100","0010","0011","0100","0100","0110","0110","0110","0101","0100","0100","0011","0011","0100","0101","0101","0101","0101","0100","0011","0100","0100","0100","0100","0101","0101","0100","0011","0100","0101","0011","0011","0010","0011","0100","0011","0101","0100","0011","0101","0101","0101","0100","0100","0101","0110","0110","0110","0101","0101","0101","0101","0100","0011","0100","0100","0011","0011","0011","0011","0011","0100","0101","0111","1001","1001","1001","1001","1000","0111","0101","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0101","0100","0100","0011","0011","0101","0101","0101","0101","0101","0110","0110","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0100","0101","0100","0011","0010","0011","0011","0011","0011","0011","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0010","0010"),
("0100","0100","0101","0011","0010","0011","0100","0100","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0110","0101","0101","0101","0100","0010","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0101","0110","0110","0100","0100","1000","0100","0010","0011","0111","0110","0011","0111","1000","1000","0111","0101","0011","0010","0010","0010","0010","0010","0001","0001","0101","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1001","1001","0111","0100","0100","0100","0100","0100","0011","0011","0011","0100","0111","1000","0111","0100","0100","0100","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0101","0100","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0011","0110","0110","0011","0010","0010","0011","0110","0101","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0011","0100","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0011","0101","0100","0100","0101","0100","0101","0011","0101","0011","0101","0011","0101","0100","0101","0100","0100","0111","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0100","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0001","0001","0001","0011","0100","0010","0011","0100","0100","0011","0011","0001","0010","0100","0100","0100","0100","0011","0011","0011","0100","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0011","0100","0011","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0100","0101","0111","1000","1001","1000","0100","0011","0011","0011","0100","0011","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0110","0111","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0101","0101","0101","0100","0100","0100","0101","0101","0100","0100","0100","0101","0101","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0101","0100","0011","0011","0011","0010","0010","0100","0100","0111","1010","1010","1000","1000","1001","1001","1001","1001","1001","0100","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0011","0100","0101","0101","0110","0101","0101","0100","0101","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010"),
("0010","0100","0101","0010","0010","0011","0011","0100","0110","0111","0111","0111","0111","0111","0101","0101","0110","0100","0101","0101","0011","0011","0100","0100","0010","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0101","0110","0110","0100","0100","1000","0100","0010","0011","0111","0110","0011","0111","1000","1000","0111","0101","0011","0011","0011","0011","0011","0011","0010","0010","0100","1000","1000","1001","1001","1000","1000","0101","1000","1000","1000","1000","1001","0111","0100","0100","0100","0100","0100","0100","0011","0011","0111","1001","1001","1001","0111","0110","0110","0101","0101","0101","0100","0100","0100","0100","0100","0011","0011","0011","0100","0011","0011","0011","0100","0101","0110","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0100","0100","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0101","0011","0001","0001","0011","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0100","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","0011","0101","0100","0100","0101","0100","0101","0011","0110","0011","0110","0011","0101","0100","0101","0100","0100","0111","0100","0100","0101","0100","0100","0100","0100","0101","0100","0101","0100","0101","0011","0101","0100","0101","0100","0101","0100","0100","0100","0100","0010","0100","0100","0100","0100","0101","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0011","0011","0100","0101","0100","0010","0001","0001","0011","0011","0010","0011","0100","0011","0011","0011","0010","0011","0100","0100","0011","0011","0011","0011","0010","0100","0110","0101","0011","0011","0010","0010","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0101","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0011","0100","0100","0101","0101","0101","0101","0100","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0011","0101","0100","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0100","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0101","0011","0100","0101","0100","0011","0101","0101","0101","0101","0110","0110","0100","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0110","0101","0100","0100","0101","0110","0101","0100","0011","0011","0011","0100","0101","0110","0110","0110","0110","0101","0011","0100","0010","0100","0101","0110","0111","0111","0110","0101","1000","1001","1010","1001","1001","1001","0100","0010","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0100","0110","0110","0110","0110","0101","0101","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010"),
("0010","0100","0101","0010","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0101","0011","0100","0101","0101","0010","0010","0100","0011","0010","0100","0100","0100","0100","0100","0101","0100","0101","0101","0100","0101","0011","0011","0100","0100","0100","0101","0101","0100","0100","0111","0011","0010","0010","0111","0110","0010","0111","1000","1000","0111","0101","0100","0011","0100","0100","0100","0101","0011","0011","0101","1000","0101","0111","1001","1000","0111","0010","0111","1000","1001","1001","1001","0111","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0110","0111","0110","0100","0110","1000","1000","1000","1000","0111","0110","0101","0101","0100","0100","0101","0100","0100","0100","0110","1001","1001","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0110","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0011","0010","0011","0011","0011","0100","0100","0011","0011","0010","0001","0001","0010","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0100","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0111","0011","0101","0100","0100","0101","0011","0101","0011","0110","0011","0110","0011","0101","0100","0101","0100","0100","0111","0101","0100","0100","0100","0100","0101","0100","0101","0100","0101","0100","0101","0011","0101","0100","0101","0100","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0011","0011","0100","0100","0100","0100","0100","0101","0100","0100","0100","0010","0011","0011","0101","0101","0010","0001","0001","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0100","0011","0011","0011","0011","0010","0101","0110","0110","0011","0011","0010","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0100","0111","0100","0100","0100","0011","0011","0100","0100","0011","0011","0100","0100","0100","0101","0100","0101","0101","0101","0100","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0101","0101","0011","0100","0100","0100","0101","0101","0100","0100","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0100","0010","0010","0010","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0011","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0100","0101","0100","0100","0100","0011","0100","0110","0100","0011","0100","0101","0110","0101","0100","0011","0010","0011","0011","0101","0101","0101","0101","0101","0101","0011","0011","0011","0011","0011","0101","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","0101","0010","0010","0011","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0101","0110","0101","0100","0100","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0011"),
("0110","0101","0100","0100","0100","0101","0101","0101","0101","0100","0100","0010","0010","0101","0100","0100","0010","0011","0100","0101","0010","0010","0100","0010","0011","0100","0011","0101","0110","0101","0111","0100","0110","0110","0100","0101","0011","0100","0100","0011","0110","0111","0100","0011","0100","0111","0101","0011","0011","0110","0110","0100","0110","0101","1000","0111","0100","0011","0010","0011","0100","0100","0101","0011","0011","0100","0111","0100","0110","1000","1000","0110","0010","0101","0111","0111","0111","1000","0110","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0101","0100","0100","0100","0100","0100","0110","0100","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0110","1000","0111","0101","0101","0100","0110","0110","0101","0011","0010","0010","0010","0010","0010","0001","0010","0010","0010","0011","0110","0110","0110","0101","0011","0011","0011","0011","0100","0011","0100","0011","0011","0010","0001","0001","0001","0011","0100","0110","0110","0100","0100","0011","0011","0011","0011","0011","0011","0011","0110","0101","0101","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0100","0100","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0010","0011","0111","0100","0101","0100","0100","0101","0100","0101","0011","0110","0011","0110","0011","0101","0100","0100","0101","0100","0111","0101","0100","0100","0101","0100","0101","0100","0101","0100","0101","0100","0101","0011","0101","0100","0101","0100","0101","0011","0011","0011","0011","0011","0101","0100","0101","0100","0100","0010","0010","0011","0100","0101","0100","0011","0101","0101","0101","0011","0010","0010","0011","0110","0101","0100","0100","0100","0101","0101","0100","0100","0100","0101","0101","0100","0101","0100","0101","0101","0101","0101","0101","0100","0100","0110","0111","0110","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0100","0101","0101","0101","0110","0101","0101","0100","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0100","0010","0010","0010","0011","0101","0110","0110","0110","0101","0101","0101","0101","0101","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0011","0011","0101","0100","0100","0011","0010","0010","0010","0011","0100","0100","0011","0011","0100","0101","0011","0010","0011","0011","0011","0100","0101","0101","0101","0101","0110","0101","0110","1000","1001","1001","0101","0011","0011","0011","0010","0010","0011","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0101","0110","0110","0110","0110","0110","0101","0011","0100","0110","0101","0110","0110","0101","0110","0110","0110"),
("0111","0101","0100","0100","0100","0100","0101","0101","0101","0110","0101","0101","0101","0101","0101","0100","0010","0011","0011","0100","0011","0100","0011","0011","0100","0100","0011","0101","0111","0111","0111","0110","0110","0110","0101","0011","0011","0011","0011","0011","0110","0101","0011","0011","0101","0110","0110","0101","0100","0100","0101","0100","0100","0011","0110","0101","0011","0011","0101","0110","0100","0100","0100","0011","0011","0100","0111","0100","0101","1000","0111","0111","0110","0110","0110","0111","0111","0111","0101","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0110","0110","0101","0011","0011","0100","0100","0011","0011","0011","0011","0010","0011","0011","0011","0100","0110","0101","0011","0011","0100","0100","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","0110","1000","1000","1000","1000","1000","1000","1000","0111","0100","0011","0100","0110","0110","0100","0011","0100","0011","0011","0011","0100","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0011","0101","0101","0101","0100","0011","0011","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0011","0101","0110","0110","0100","0011","0011","0010","0011","0010","0011","0011","0101","0110","0101","0101","0101","0011","0010","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0011","0100","0101","0100","0011","0011","0011","0100","0010","0010","0010","0011","0011","0011","0011","0011","0011","0111","0100","0101","0101","0100","0101","0100","0110","0011","0110","0011","0110","0011","0101","0100","0101","0101","0100","0111","0101","0100","0101","0101","0101","0101","0100","0101","0100","0110","0100","0101","0011","0101","0100","0101","0100","0101","0011","0010","0011","0011","0010","0100","0100","0100","0011","0011","0010","0010","0011","0100","0011","0011","0011","0011","0100","0100","0011","0011","0010","0011","0100","0100","0100","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0100","0100","0100","0100","0101","0100","0100","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0101","0100","0011","0100","0100","0010","0010","0010","0011","0101","0101","0110","0110","0101","0101","0110","0111","0101","0110","0101","0100","0100","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0110","0110","0110","0100","0010","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0010","0011","0010","0011","0100","0101","0100","0101","0110","0100","0011","0100","0101","0011","0011","0011","0100","0011","0011","0011","0010","0010","0010","0011","0100","0010","0010","0010","0100","0100","0011","0010","0010","0011","0011","0011","0010","0010","0100","0011","0001","0010","0110","1001","1001","1001","0100","0010","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0011","0100","0110","0111","0111","0111","0111","0110","0111","0110","0010","0010","0001","0101","0110","0110","0110","0110","0110","0110","0110"),
("0011","0010","0010","0010","0010","0010","0010","0011","0100","0110","0111","0111","0111","0110","0100","0011","0010","0010","0011","0100","0101","0101","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0011","0100","0011","0011","0101","0101","0100","0101","0100","0100","0101","0101","0101","0101","0110","0110","0110","0110","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0111","1000","0101","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0010","0100","0110","0100","0011","0010","0011","0011","0101","1000","1001","0111","0110","0101","0101","0101","0101","0110","0100","0100","0110","0100","0100","0101","0101","0100","0101","0100","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0011","0011","0011","0010","0010","0010","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0011","0100","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0110","0110","0101","0101","0101","0100","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","0100","0101","0100","0100","0101","0011","0110","0011","0110","0011","0110","0011","0101","0100","0100","0101","0011","0111","0101","0100","0101","0101","0101","0101","0100","0101","0100","0101","0100","0101","0100","0101","0100","0101","0100","0101","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0101","0100","0100","0100","0101","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0100","0100","0011","0011","0011","0100","0010","0010","0010","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0110","0100","0100","0100","0011","0010","0010","0100","0100","0100","0100","0011","0011","0011","0011","0101","0101","0101","0101","0101","0100","0010","0010","0010","0010","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0110","1000","0100","0010","0011","0100","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0100","0100","0011","0011","0011","0111","0101","0010","0011","0111","1000","1000","1000","0101","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0011","0010","0010","0010","0010","0010","0100","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0100","0010","0010","0001","0011","0110","0110","0110","0110","0110","0110","0110"),
("0010","0001","0011","0011","0010","0010","0011","0100","0011","0100","0101","0011","0010","0100","0100","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0011","0010","0010","0001","0010","0010","0010","0010","0100","0100","0011","0011","0011","0011","0100","0100","0011","0100","0110","0101","0101","0111","0011","0101","0110","0101","0011","0010","0011","0100","0100","0100","0100","0011","0010","0010","0010","0110","0110","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0100","0011","0010","0010","0011","0011","0010","0100","0101","0100","0011","0100","0100","0100","0100","0100","0011","0100","0101","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","0101","0110","0110","0101","0101","0100","0100","0100","0100","0011","0100","0100","0110","0111","0111","0111","0111","0111","0111","0111","0110","0101","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0111","0110","0111","0111","0111","0111","0110","0111","0110","0111","0110","0111","0110","0111","0111","0111","0111","0110","0111","0110","0101","0110","0101","0110","0101","0110","0110","0101","0101","0101","0110","0101","0110","0101","0110","0100","0101","0100","0100","0100","0100","0100","0101","0101","0101","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0010","0011","0010","0011","0100","0100","0100","0110","0101","0100","0101","0100","0100","0101","0101","0100","0100","0011","0010","0010","0011","0100","0100","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0101","0111","0100","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0010","0010","0011","0111","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0110","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0011","0100","0010","0010","0100","0100","0011","0010","0010","0010","0100","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0011","0011","0010","0010","0010","0100","0110","0110","0110","0110","0110","0110"),
("0101","0100","0100","0010","0011","0101","0101","0110","0101","0101","0110","0011","0001","0101","0101","0011","0011","0010","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0110","0101","0100","0100","0100","0100","0100","0101","0101","0101","0100","0101","0100","0011","0011","0010","0001","0001","0011","0011","0011","0011","0011","0010","0001","0010","0010","0011","0011","0011","0011","0110","0110","0101","0111","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0101","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0011","0010","0010","0011","0011","0011","0011","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0110","0101","0110","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0111","1001","1001","1000","1000","1000","1000","1000","1000","0110","0011","0100","0010","0010","0011","0100","0010","0010","0010","0010","0011","0011","0010","0111","1001","1001","1001","1001","1000","1001","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1000","1000","0101","0100","0101","0100","0100","0100","0100","0101","0100","0101","0100","0101","0100","0101","0100","0101","0100","0101","0100","0100","0100","0100","0100","0101","0101","0101","0011","0011","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0101","0101","0101","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0011","0100","0101","0100","0011","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0011","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0011","0011","0100","0011","0110","0111","0110","0110","0101","0101","0110","0011","0011","0010","0010","0010","0011","0100","0100","0100","0100","0011","0100","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0111","0101","0101","0011","0100","0100","0101","0100","0011","0011","0100","0101","0101","0101","0101","0110","0101","0011","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0010","0010","0011","1001","1010","1010","1010","1010","1010","1010","1010","1001","1001","1000","1000","1000","1000","0111","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0011","0011","0010","0010","0010","0010","0010","0011","0100","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0100","0010","0010","0001","0010","0010","0011","0110","0111","0111","0110","0111","0110"),
("0101","0101","0100","0010","0011","0101","0101","0101","0110","0111","0110","0110","0110","0110","0100","0100","0100","0011","0100","0101","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0110","0110","0101","0110","0101","0110","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0100","0011","0010","0010","0010","0011","0100","0011","0100","0011","0011","0001","0010","0011","0011","0011","0011","0011","0101","0111","1000","1000","0101","0100","0011","0011","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0100","0100","0101","0101","0101","0100","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0001","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0111","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0111","1000","1000","1000","1000","1000","1000","1000","1000","0110","0011","0100","0010","0010","0011","0100","0010","0010","0010","0010","0100","0011","0010","0111","1000","1001","1001","1000","1001","1001","1000","1001","1001","1001","1000","1001","1000","1000","1000","1001","1000","0111","0101","0100","0101","0100","0101","0101","0100","0101","0100","0101","0100","0101","0100","0101","0100","0101","0100","0101","0100","0011","0011","0011","0010","0011","0011","0011","0010","0011","0011","0011","0001","0011","0010","0010","0010","0001","0001","0010","0100","0001","0011","0100","0101","0101","0101","0101","0101","0101","0110","0110","0110","0101","0101","0110","0101","0100","0100","0101","0101","0100","0100","0100","0101","0100","0100","0101","0101","0100","0100","0100","0011","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0011","0010","0001","0010","0010","0001","0001","0010","0010","0001","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0001","0010","0010","0010","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","0011","0011","0011","0010","0010","0111","1000","0110","0101","0101","0100","0100","0011","0010","0010","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0101","0111","1000","0111","0111","1000","0111","0111","0111","0111","0101","0100","0100","0110","0101","0101","0011","0011","0011","0100","0101","0101","0101","0100","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0011","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","0111","0110","0110","1000","0111","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0001","0010","0010","0010","0100","0110","0111","0111","0110","0110","0110","0100","0110","0111","0111","0111","0110","0111","0111","0111","0110","0100","0011","0011","0011","0010","0100","0111","0110","0110","0111","0110","0111"),
("0010","0001","0001","0011","0011","0010","0011","0100","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0101","0110","0110","0110","0110","0110","0110","0101","0101","0101","0100","0100","0100","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0101","0100","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0011","0100","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0101","0100","0100","0011","0100","0100","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0011","0100","0111","1000","1000","1000","1000","1000","1000","1000","1000","0101","0010","0100","0001","0001","0100","0100","0001","0001","0001","0010","0100","0011","0010","0111","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","0111","0101","0100","0101","0100","0100","0101","0100","0101","0100","0101","0100","0101","0011","0101","0100","0101","0100","0101","0011","0011","0011","0011","0010","0100","0011","0011","0010","0011","0011","0011","0010","0011","0010","0011","0011","0010","0010","0010","0100","0010","0100","0100","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0101","0101","0101","0101","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0001","0011","0010","0001","0010","0011","0100","0100","0100","0101","0101","0110","0110","0101","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0110","0110","0100","0011","0100","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0100","0101","0100","0101","0101","0101","1000","1000","1000","0110","0101","0110","0101","0011","0101","0101","0100","0100","0011","0010","0100","0100","0011","0100","0011","0011","0011","0100","0011","0010","0010","0010","0010","0010","0011","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1000","1000","1000","1001","1000","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0010","0011","0100","0100","0101","0110","0111","0111","0110","0110","0110","0100","0110","0111","0111","0111","0111","0111","0111","0111","0101","0011","0010","0010","0010","0010","0011","0110","0100","0100","0110","0100","0011"),
("0011","0001","0001","0100","0011","0010","0100","0101","0100","0010","0010","0001","0010","0010","0011","0100","0100","0011","0100","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0110","0110","0101","0101","0100","0100","0100","0011","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0100","0101","0100","0011","0100","0100","0100","0100","0100","0100","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0011","0011","0100","0110","1000","1000","1000","1000","1000","1001","1000","1000","0101","0010","0100","0001","0010","0100","0100","0001","0001","0001","0010","0100","0011","0010","0111","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1000","1000","1000","1001","1000","1000","1000","0111","0101","0100","0101","0101","0100","0101","0100","0101","0100","0101","0101","0110","0011","0101","0100","0101","0100","0101","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0101","0101","0110","0110","0110","0111","0110","0110","0110","0101","0101","0110","0110","0101","0101","0101","0101","0110","0110","0101","0101","0110","0101","0100","0100","0100","0101","0110","0110","0110","0110","0110","0101","0100","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0101","0111","0111","0101","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0010","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0100","0100","0101","0100","0100","0101","1000","1000","1000","0101","0101","0110","0100","0010","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0100","0011","0011","0010","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","1001","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1000","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0011","0011","0010","0010","0010","0010","0011","0100","0100","0101","0101","0101","0110","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0100","0011","0010","0010","0010","0010","0110","0110","0110","0110","0100","0010"),
("0101","0100","0011","0010","0100","0101","0101","0101","0110","0101","0011","0011","0100","0100","0011","0011","0011","0100","0100","0101","0101","0101","0101","0101","0110","0101","0101","0101","0100","0100","0100","0110","0110","0110","0111","0110","0101","0100","0100","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0100","0100","0100","0011","0010","0010","0100","0011","0011","0011","0011","0010","0010","0010","0011","0011","0100","0011","0011","0100","0100","0100","0101","0100","0100","0011","0011","0011","0100","0011","0100","0011","0011","0011","0100","0100","0110","0111","0110","0011","0011","0011","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0110","0101","0101","0100","0101","0101","0100","0101","0101","0101","0100","0100","0011","0100","0100","0110","1000","1000","1000","1000","1000","1000","1000","1000","0110","0010","0100","0010","0010","0100","0100","0010","0010","0010","0011","0100","0010","0010","0111","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","0101","0100","0101","0101","0100","0101","0100","0101","0100","0101","0101","0101","0011","0101","0100","0110","0100","0101","0101","0100","0100","0100","0100","0101","0101","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0101","0101","0110","0110","0110","0111","0110","0100","0010","0010","0011","0101","0110","0111","0110","0110","0110","0101","0101","0101","0110","0100","0100","0100","0101","0101","0101","0110","0110","0101","0011","0001","0001","0010","0100","0110","0110","0111","0110","0110","0101","0011","0100","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0011","0010","0001","0010","0010","0010","0010","0010","0001","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0100","0100","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0100","0100","0101","0110","0111","1000","1000","0110","0101","0110","0100","0011","0010","0010","0011","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0100","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","1001","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1010","1001","0110","0011","0010","0011","0100","0100","0011","0011","0010","0010","0100","0011","0010","0010","0010","0010","0010","0011","0101","0101","0101","0011","0010","0010","0010","0010","0010","0011","0101","0101","0101","0011","0010","0010","0010","0010","0001","0011","0101","0100","0011","0010","0010","0010","0100","0010","0010","0010","0010","0010","0010","0010","0100","0011","0010","0010","0010","0011","0011","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0100","0100","0100","0011","0010","0010","0011","0010","0011","0100","0101","0110","0101","0101","0110","0110","0110","0110","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0100","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0010"),
("0101","0100","0011","0010","0011","0100","0100","0100","0101","0100","0100","0110","0110","0110","0100","0011","0100","0100","0100","0101","0101","0101","0101","0101","0101","0011","0010","0011","0011","0011","0011","0101","0101","0110","0110","0110","0110","0101","0101","0110","0110","0111","0110","0111","0111","0111","0111","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0100","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","0110","0011","0011","0011","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0101","0101","0101","0101","0110","0110","0101","0110","0110","0110","0100","0100","0011","0100","0100","0110","1000","1000","1000","1000","1000","1000","1000","1000","0110","0101","0101","0100","0101","0101","0101","0100","0101","0100","0100","0011","0010","0010","0110","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","0110","0101","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0101","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0010","0011","0011","0011","0010","0010","0010","0011","0011","0010","0011","0011","0011","0010","0100","0101","0101","0100","0100","0100","0110","0110","0110","0110","0111","0100","0010","0010","0001","0001","0010","0101","0111","0111","0111","0110","0101","0101","0101","0101","0100","0100","0101","0110","0101","0101","0101","0110","0011","0001","0000","0001","0001","0010","0101","0110","0110","0110","0110","0100","0011","0100","0101","0010","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0011","0011","0101","0110","0111","1000","1000","1000","0100","0100","0101","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0011","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0011","0010","0011","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","0101","0010","0001","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0010","0011","0100","0011","0011","0011","0011","0011","0100","0100","0100","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0101","0101","0101","0101","0011","0011","0100","0011","0101","0101","0100","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0100","1010","1011","1011","1011","1000","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0101","0101","0101","0110","0110","0110","0110","0110","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001"),
("0010","0001","0001","0010","0010","0001","0001","0010","0011","0100","0101","0101","0110","0110","0101","0100","0100","0011","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0110","0101","0101","0110","0110","0110","0110","0101","0110","0111","0111","0110","0111","0111","0111","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0111","0111","0110","0110","0101","0100","0100","0011","0010","0010","0011","0011","0011","0011","0010","0010","0001","0010","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0110","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0100","0100","0110","1000","1000","1000","1001","1001","1001","1000","1000","0110","0011","0100","0011","0100","0011","0100","0011","0100","0011","0011","0010","0010","0010","0110","0111","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","0110","0100","0101","0100","0101","0100","0100","0100","0100","0101","0100","0101","0100","0101","0100","0101","0100","0101","0100","0011","0011","0011","0010","0100","0011","0011","0010","0011","0011","0011","0001","0001","0001","0011","0100","0001","0011","0010","0100","0010","0011","0101","0101","0101","0100","0100","0101","0110","0110","0110","0110","0011","0010","0001","0001","0001","0001","0011","0111","0110","0110","0110","0110","0101","0101","0110","0100","0101","0110","0110","0101","0101","0101","0100","0001","0001","0001","0000","0001","0010","0100","0110","0110","0110","0101","0101","0100","0100","0101","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0100","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0101","0110","1000","1000","0111","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0101","0101","0100","0011","0010","0010","0010","0010","0011","0010","0100","0110","0110","0100","0010","0010","0010","0010","0010","0011","0011","0011","0101","0011","0010","0010","0010","0011","0101","0100","0010","0011","0110","0110","0110","0110","0100","0010","0010","0011","0110","0111","0101","0010","0010","0010","0010","0010","0101","0110","0101","0100","0101","0100","0101","0101","0101","0101","0101","0100","0100","0100","0101","1000","0111","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0110","0110","0101","0101","0100","0010","0011","0011","0011","0010","0001","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0001"),
("0100","0010","0010","0011","0011","0011","0011","0100","0011","0100","0101","0011","0011","0101","0101","0011","0010","0010","0001","0010","0011","0100","0100","0101","0110","0110","0110","0101","0011","0101","0101","0101","0101","0101","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0101","0100","0100","0011","0010","0011","0100","0100","0100","0100","0011","0011","0010","0010","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0101","0101","0110","0110","0110","0111","0110","0110","0110","0110","0110","0101","0100","0100","0100","0100","0111","1000","1000","1000","1000","1000","1000","1000","1000","0110","0011","0100","0011","0100","0011","0100","0011","0100","0011","0011","0011","0010","0010","0110","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0110","0100","0101","0100","0101","0100","0100","0101","0100","0101","0100","0101","0100","0101","0100","0110","0100","0110","0101","0101","0101","0101","0101","0110","0110","0110","0111","0111","0110","0111","0111","0111","0111","0101","0101","1000","1001","1001","1001","1001","1001","1010","1000","0110","0100","0100","0101","0110","0110","0110","0101","0011","0011","0001","0001","0010","0010","0010","0110","0110","0110","0110","0110","0101","0101","0101","0100","0101","0110","0110","0101","0101","0110","0100","0001","0001","0001","0001","0001","0010","0011","0101","0110","0110","0101","0100","0100","0101","0110","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0001","0001","0010","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0111","1000","0111","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0010","0101","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0011","0011","0100","0101","0110","0111","1000","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","0110","0111","0111","0110","0110","0110","0110","0110","0111","0110","0101","0110","0110","0110","0101","0110","0100","0100","0100","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0110","1100","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0110","0110","0110","0100","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0101","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0010","0001","0001","0001","0001","0010","0011","0011","0011","0100","0100","0100","0100","0011","0100","0101","0101","0101","0100","0101","0110","0110","0101","0101","0110","0110","0101","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","0101","0110","0111","0110","0110","0110","0110","0110","0111","0111","0110","0110","0100","0100","0100","0100","0110","1000","1000","1000","1000","1000","1000","1000","1000","0110","0010","0100","0011","0100","0100","0100","0011","0100","0011","0011","0011","0010","0010","0110","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0110","0100","0101","0101","0101","0101","0100","0101","0100","0110","0101","0110","0110","0111","0111","1000","1000","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1000","0110","1010","1010","1010","1001","1000","1000","1000","0111","0110","0100","0100","0100","0101","0110","0110","0101","0011","0011","0001","0001","0010","0010","0010","0101","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0110","0110","0101","0110","0100","0001","0001","0001","0000","0001","0011","0011","0101","0110","0110","0101","0100","0100","0101","0101","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0110","0111","1000","0101","0101","0101","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0010","0011","0010","0010","0011","0011","0010","0011","0010","0100","0101","0100","0011","0010","0010","0100","1010","1011","1011","1010","1010","1000","0111","0110","0110","1001","1010","1010","1010","1010","1000","0011","0101","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0110","0101","0101","0110","0011","0010","0010","0100","0111","0111","0110","0110","0111","0110","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1001","0111","0110","0101","0101","0110","0111","0110","0011","0011","0011","0011","0011","0011","0010","0011","0010","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010"),
("0101","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0111","0110","0011","0010","0001","0010","0010","0010","0001","0001","0001","0011","0011","0010","0011","0011","0011","0010","0010","0011","0101","0110","0101","0101","0110","0111","0110","0101","0110","0110","0101","0101","0101","0110","0110","0110","0111","1000","1001","1001","1001","0111","0101","0101","0110","0101","0101","0101","0101","0100","0100","0100","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0110","0110","0111","0111","0110","0110","0110","0111","0111","0111","0110","0110","0101","0100","0100","0100","0110","1000","1000","1000","1000","1000","1001","1000","0110","0110","0011","0100","0100","0100","0100","0100","0011","0100","0100","0011","0100","0010","0010","0111","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0110","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0011","0011","0011","0011","0101","0101","0100","0011","0101","0110","0110","0110","0101","0100","0011","0001","0001","0010","0010","0010","0101","0110","0110","0101","0101","0100","0100","0101","0101","0100","0101","0101","0110","0110","0110","0011","0001","0010","0010","0001","0010","0100","0100","0110","0110","0110","0101","0100","0011","0101","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0001","0010","0010","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0101","0110","0111","0111","0110","0101","0011","0010","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0101","0110","0110","0110","0110","0110","0110","0101","0101","0110","1010","1010","1010","1011","1001","0100","0011","0011","0011","0110","1010","1010","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","0110","0110","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","0111","0111","0101","0011","0010","0010","0010","0011","0101","0110","0011","0011","0101","0100","0100","0111","0111","0111","0111","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0100","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0001","0001","0010","0001","0001","0001","0010","0011","0011","0011","0011","0010","0010"),
("0110","0011","0010","0101","0100","0010","0011","0101","0100","0100","0101","0101","0100","0010","0001","0010","0010","0010","0010","0001","0001","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0100","0110","0110","0110","0110","0110","0110","0100","0100","0101","0101","0110","0110","0110","0110","0110","0110","0111","1000","1000","0111","0110","0110","0110","0101","0101","0101","0101","0100","0100","0100","0100","0011","0010","0010","0100","0100","0011","0100","0011","0011","0010","0010","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0011","0011","0100","0101","0100","0100","0100","0010","0011","0011","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0011","0011","0100","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0100","0100","0100","0101","0101","0110","0110","0110","1000","0111","0110","0110","0010","0100","0100","0100","0011","0100","0011","0100","0011","0011","0011","0010","0010","0110","1000","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0110","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0101","0101","0100","0101","0101","0101","0100","0011","0101","0110","0110","0111","0110","0101","0100","0010","0010","0011","0011","0011","0110","0110","0110","0101","0101","0100","0100","0101","0100","0100","0101","0101","0101","0110","0110","0100","0010","0010","0010","0001","0011","0100","0100","0110","0110","0110","0101","0100","0011","0101","0101","0010","0001","0001","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0001","0010","0010","0010","0010","0010","0001","0001","0010","0001","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0101","0101","0111","0111","0110","0110","0110","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0110","0111","0111","1000","1000","0111","1000","0111","0111","0111","1010","1011","1011","1001","0011","0010","0010","0010","0010","0100","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0100","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0110","0101","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0101","0110","1000","1000","1000","1000","1000","0111","0010","0010","0010","0011","0111","0110","0111","0101","0010","0011","0010","0010","0010","0010","0100","1000","1000","1000","1000","0111","0011","0101","1000","0111","0110","0100","0010","0010","0010","0010","0010","0010","0101","0100","0010","0010","0011","0011","0011","0010","0010","0001","0001","0010","0010","0010","0001","0001","0100","0100","0011","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010"),
("0110","0100","0011","0101","0100","0011","0100","0100","0100","0100","0101","0100","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0011","0011","0010","0010","0010","0010","0010","0010","0010","0100","0101","0101","0101","0110","0110","0101","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0100","0101","0101","0101","0101","0101","0100","0101","0011","0010","0011","0011","0100","0011","0010","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0101","0101","0100","0011","0011","0100","0011","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0011","0100","0101","0110","0110","0110","0110","0110","0101","0100","0101","0101","0101","0101","0101","0100","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0101","0100","0101","0100","0100","0100","0100","0011","0011","0011","0010","0010","0110","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0111","0101","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0110","0101","0110","0110","0100","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0100","0011","0011","0111","1000","1000","1000","1000","0111","1000","0110","0101","0101","0100","0101","0110","0110","0111","0111","0101","0110","0011","0001","0011","0010","0011","0111","0111","0110","0101","0101","0101","0100","0101","0100","0100","0110","0110","0110","0101","0110","0101","0010","0001","0010","0001","0100","0101","0101","0110","0110","0110","0101","0100","0100","0101","0101","0010","0001","0001","0001","0010","0001","0001","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0011","0010","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0101","0101","0101","0110","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0100","0011","0011","0010","0010","0010","0011","0101","0100","0110","0110","0110","0110","0110","0111","0110","0111","0110","1010","1010","1001","1000","0100","0010","0010","0011","0100","0110","1000","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","0011","0001","0001","0100","1000","0110","0111","0110","0010","0010","0010","0010","0010","0001","0100","1000","1000","1000","1001","1000","0010","0100","1000","0111","0110","0101","0100","0011","0010","0010","0001","0001","0011","0011","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0011","0010","0010","0100","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010"),
("0101","0100","0100","0101","0101","0100","0011","0100","0011","0100","0101","0101","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0011","0100","0011","0010","0010","0011","0010","0010","0010","0011","0100","0100","0100","0101","0101","0101","0100","0011","0100","0100","0011","0100","0100","0100","0101","0101","0100","0100","0011","0100","0101","0101","0100","0100","0101","0100","0101","0101","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0100","0011","0101","0111","0111","0110","0110","0110","0101","0110","0110","0101","0101","0101","0100","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0101","0110","0110","0111","0110","0111","0111","0111","0110","0110","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0010","0011","0010","0011","0010","0011","0010","0010","0010","0110","1000","1000","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","0111","0101","0110","0101","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0010","0101","0110","0110","0110","0110","0110","0110","0101","0101","0101","0100","0100","0101","0100","0011","1000","1001","1001","1001","1001","1010","1010","0111","0101","0101","0100","0101","0110","0111","0111","0111","0110","0110","0110","0011","0010","0010","0101","0111","0111","0110","0110","0110","0101","0101","0101","0100","0101","0110","0111","0110","0101","0110","0101","0011","0010","0011","0100","0101","0101","0110","0110","0110","0110","0110","0100","0100","0101","0101","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0011","0010","0011","0011","0011","0010","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0101","0110","0110","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0110","0111","0111","0111","0111","0111","0110","0011","0011","0011","0010","0001","0100","0101","0100","0110","0101","0100","0100","0100","0100","0011","0010","0011","1001","0111","0100","0100","0100","0101","0101","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0101","0101","0101","0101","0101","0011","0011","0011","0011","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0101","0101","0101","0101","0101","0011","0100","0101","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0010","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001"),
("0100","0100","0011","0100","0101","0100","0011","0100","0011","0100","0101","0100","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0100","0100","0100","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0110","0110","0111","0101","0010","0011","0100","0100","0101","0110","0110","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0110","0101","0110","0110","0110","0111","0111","0110","0111","0111","0111","0110","0110","0110","0110","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0011","0010","0011","0010","0010","0001","0110","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0110","0111","1001","1001","0111","0101","0110","0100","0101","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0100","0101","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","1000","0111","0111","0111","0111","0111","0111","0110","0101","0101","0100","0101","0110","0110","0110","0111","0111","0111","0111","0111","0110","0110","0110","0111","0110","0110","0110","0110","0101","0100","0101","0101","0101","0110","0110","0110","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0100","0101","0101","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0101","0111","1000","1000","1000","1000","1001","1001","1001","1000","0111","0101","0011","0010","0010","0100","0101","0101","0101","0101","0011","0010","0011","0011","0010","0010","0010","1000","0111","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0100","0100","0011","0010","0011","0101","0101","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0011","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0010","0011","0010","0010","0001","0001"),
("0101","0100","0100","0100","0100","0011","0011","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0011","0010","0011","0011","0011","0010","0010","0011","0010","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0110","0110","0101","0110","0101","0100","0100","0101","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0100","0110","0111","0110","0110","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0001","0110","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0110","0101","1000","1001","0111","0100","0110","0101","0110","0101","0101","0101","0111","0110","0110","0110","0110","0101","0101","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","1000","0101","0100","0011","0011","0111","1000","0110","0101","0100","0100","0101","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0110","0110","0101","0100","0101","0101","0100","0110","0110","0101","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0101","0101","0010","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0010","0011","0110","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1001","1000","1001","1000","0110","0110","0111","0111","0111","0111","0111","0100","0010","0011","0101","0100","0101","0101","0110","0110","0110","0101","0100","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0100","0011","0001","0001","0010","0100","0100","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0010","0010","0011","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0001"),
("0101","0100","0011","0011","0100","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0001","0001","0010","0001","0010","0011","0011","0010","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0100","0011","0100","0100","0011","0011","0011","0110","1000","1000","1001","0111","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","0110","0110","0110","0110","0110","0111","0111","0110","0011","0010","0100","0110","0110","0110","0111","0111","0110","0101","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0001","0110","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0110","0100","0111","1000","0111","0100","0110","0101","0110","0101","0101","0101","0110","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","1000","0101","0011","0010","0010","0111","1000","0111","0101","0101","0100","0101","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0101","0101","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0011","0011","0010","0010","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0100","0110","1000","1001","1001","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1000","1001","1000","1001","1000","1000","1000","1000","1000","1001","0100","0010","0100","0110","0111","1000","1000","0111","0111","1000","0111","0110","0111","0110","0100","0100","0100","0100","0100","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0010","0001","0010","0011","0011","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010"),
("0101","0100","0011","0011","0100","0011","0011","0011","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0010","0010","0011","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0011","0110","1000","1000","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0101","0110","0111","0110","0111","0111","0110","0110","0101","0100","0011","0100","0110","0111","0111","0111","0111","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0110","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0110","0011","0111","1001","0111","0110","0111","0110","0110","0101","0100","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0101","0101","0100","0100","0101","0101","0110","0101","1000","0110","0100","0011","0011","0111","1000","0111","0110","0101","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0101","0110","0101","0101","0111","0111","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0101","0101","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0001","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0100","0110","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0110","0100","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0101","0111","1001","1001","1001","1000","1001","1000","0111","0101","0111","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","0101","0100","0101","0111","1000","0111","0111","0111","0111","0110","1000","0101","0101","0101","0100","0011","0011","0011","0011","0100","0100","0011","0011","0011","0100","0100","0100","0011","0011","0100","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0010","0001","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010"),
("0101","0011","0010","0011","0011","0011","0011","0100","0011","0010","0010","0011","0011","0010","0010","0011","0010","0010","0010","0001","0001","0001","0010","0001","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0011","0011","0010","0001","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0101","0100","0011","0011","0100","0101","0101","0100","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0110","0100","0101","0110","0111","0111","0111","0110","0110","0110","0101","0100","0101","0111","0111","0111","0110","0111","0110","0110","0110","0101","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0110","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","0111","0111","1000","0110","0100","0110","0111","0111","0111","0111","0111","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0101","0110","0101","0101","0101","0101","0101","0110","0110","0110","0101","0100","0101","0110","0111","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0110","0110","0110","0101","0110","0101","0101","0111","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0101","0110","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0101","0101","0011","0010","0010","0010","0011","0011","0011","0100","0100","0100","0100","0101","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0110","0100","0010","0010","0100","0100","0100","0011","0011","0011","0101","0110","1000","1001","1001","1001","1001","1000","1001","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","0111","1000","0111","0101","0110","0111","0111","0111","0111","0111","0110","0111","0111","0101","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0100","0100","0100","0100","0100","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0011","0010","0011","0100","0011","0011","0011","0100","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0010","0011","0011","0011","0011","0011","0010","0010","0010","0001","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0011","0011","0100","0100","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0110","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0101","0011","0100","0110","0111","0111","0111","0110","0110","0101","0100","0101","0101","0110","0110","0111","1001","0111","0110","0110","0110","0101","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0100","0111","0111","0111","0111","1000","0111","1000","1000","1000","1000","0111","1000","0111","0110","0110","0111","0101","0100","0100","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0100","0100","0011","0111","1010","1000","0011","0011","0011","0010","0010","0011","0101","0110","0101","0100","0101","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0110","0101","0101","0101","0101","0111","0111","0110","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0101","0100","0101","0110","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0011","0100","0100","0100","0100","0101","0110","0110","0110","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0110","0101","0100","0101","0100","0100","0100","0100","0100","0101","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0110","0110","0110","0110","0110","0110","0110","0111","0111","0101","0110","0111","0111","0110","0101","0011","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","1000","1000","1000","0110","0100","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0010"),
("0100","0101","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0010","0011","0011","0011","0011","0010","0010","0010","0010","0001","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0010","0010","0011","0011","0010","0001","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0011","0010","0001","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0011","0011","0100","0110","0111","0110","0110","0110","0110","0101","0100","0100","0101","0110","0110","0110","1001","0101","0110","0110","0110","0101","0100","0110","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0101","0110","0101","0100","0100","0110","1010","1001","0110","0011","0011","0100","0011","0011","0101","1010","1010","0111","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","1001","1010","1001","1001","1011","1010","0101","0011","0010","0010","0010","0111","1000","0110","0101","0100","0110","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0110","0110","0101","0110","0110","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0110","0110","0110","0110","0111","0111","0111","0111","0101","0101","0110","0111","0101","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0110","0111","0111","0111","0110","0111","0110","0011","0011","0100","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","0101","0101","0110","0101","0101","0101","0101","0100","0100","0011","0100","0100","0011","0101","0110","0110","0110","0101","0101","0101","0101","0110","0111","0110","0110","0100","0100","0100","0100","0100","0100","0110","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0100","0100","0100","0100","0100","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0100","0100","0110","1000","1000","0110","0110","0110","0111","1000","0110","0100","0011","0011","0011","0010","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0100","0011","0010","0011","0010","0010","0010","0010","0010","0011","0010","0011","0010"),
("0101","0101","0101","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0001","0010","0001","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0011","0010","0010","0011","0010","0011","0100","0100","0100","0100","0101","0011","0010","0010","0010","0011","0011","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0100","0010","0110","0011","0101","0101","0101","0100","0101","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1010","1010","1010","1010","1000","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0101","0110","0110","0111","1000","1000","0111","0110","0100","0100","0100","0011","0011","0011","1000","1100","1100","0111","0011","0011","0011","0011","0011","0101","1100","1100","1000","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","1100","1100","1011","0110","1000","1010","0111","0101","0100","0100","0100","1000","1001","0111","0110","0101","0110","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","0111","0110","0111","0111","0111","1000","1001","1001","0111","0111","0111","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0010","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0111","0111","0111","0111","0111","0110","0111","0110","0011","0011","0100","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0100","0011","0011","0110","0011","0011","0110","0100","0011","0101","0101","0011","0100","0101","0011","0100","0110","0011","0100","0110","0011","0100","0110","0100","0011","0100","0100","0011","0011","0011","0100","0101","0110","0110","0110","0111","0100","0101","0110","0110","0110","0110","0100","0100","0100","0100","0100","0100","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0011","0100","0100","0100","0100","0100","0100","0100","0011","0101","0100","0011","0100","0100","0100","0100","0100","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0100","0101","0111","1000","0111","0101","0101","1000","1011","1001","0101","0110","1000","1000","0110","0100","0100","0100","0011","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0100","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0010","0010","0010"),
("0101","0101","0101","0101","0100","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0001","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0100","0111","0111","0111","0111","0111","1000","0111","0111","1000","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1000","0111","0111","0110","0101","0100","0100","0100","0011","0011","0011","0100","0100","0100","0110","0110","0100","0101","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0111","1000","0110","0100","0110","0101","0110","1001","0110","0110","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0011","0011","0011","0011","0011","0100","0100","0011","0011","0100","0100","0011","0011","0100","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0101","0100","0100","0011","0011","0100","0101","0101","0101","0101","0101","0101","0110","0110","0110","0100","0010","0100","0011","0101","0110","0110","0100","0110","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","0101","0100","0100","0100","0101","0011","0101","0110","0101","0101","0101","0101","0101","0110","0111","0111","0111","0110","0100","0011","0011","0011","0011","0011","0111","1010","1010","0111","0100","0100","0100","0100","0100","0101","1010","1010","1000","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0101","1010","1011","1010","0101","0100","1001","0110","0100","0101","0100","0100","0110","0100","0011","0011","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0110","0111","0111","0111","0111","0110","0111","0111","0110","0011","0010","0100","0110","0111","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0100","0011","0011","0110","0101","0101","0110","0100","0100","0101","0101","0011","0100","0101","0100","0100","0100","0011","0100","0110","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0110","0111","0111","0101","0101","0110","0101","0111","0101","0101","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0111","1000","0111","0101","0101","0111","1000","1001","1001","1000","1000","0111","0110","0110","1000","1000","0110","0100","0100","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010"),
("0101","0101","0101","0101","0110","0100","0011","0010","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0100","0101","0110","0111","0111","0111","1000","1001","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1001","1001","1000","1000","0111","0110","0110","0101","0110","0101","0100","0110","0110","0110","0110","0111","0111","0110","0111","1000","1000","1000","1000","1000","1000","1001","0111","0110","0110","0110","0111","1001","1001","0111","0101","0100","0100","0110","0111","0111","0111","0110","0110","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0101","0100","0101","0100","0110","0110","0110","0110","0110","0101","0101","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0101","0101","0101","0101","0110","0110","0101","0110","0110","0101","0110","0110","0110","0110","0101","0101","0100","0100","0100","0100","0101","0101","0011","0011","0011","0101","0110","1000","0110","0110","0110","0110","0110","0110","0110","0101","0011","0010","0011","0101","0110","0101","0100","0111","1010","1000","1010","1001","1010","1000","1000","1010","0111","1010","0111","0111","1001","0101","1001","0110","0111","1001","0101","1000","0101","0100","0100","0101","0101","0100","0101","0100","0100","0100","0100","0101","0011","0110","0111","0111","0110","0100","0011","0010","0011","0011","0011","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0101","0101","0100","0100","0100","0100","0110","0101","0101","0100","0011","0011","0100","0101","0110","0110","0101","0110","0110","0101","0101","0101","0101","0110","0110","0110","0100","0100","0100","0010","0011","0100","0011","0100","0100","0100","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0100","0011","0100","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0111","0111","0111","0111","0111","0111","0110","0011","0010","0100","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0100","0110","0111","0110","0111","0111","0110","0110","0111","0110","0110","0111","0110","0110","0101","0110","0101","0011","0110","0110","0111","0110","0101","0110","0101","0101","0100","0011","0100","0100","0101","0110","0110","0100","0101","0101","0110","0101","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0011","0011","0011","0100","0100","0001","0010","0011","0011","0011","0011","0011","0011","0011","0100","0101","0111","1000","0111","0101","0101","0110","0111","1000","1000","1000","1000","1000","0110","1001","0111","0110","0110","0110","1000","1000","0110","0100","0100","0011","0010","0010","0010","0011","0011","0011","0011","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0010","0010","0010"),
("0110","0110","0110","0110","0110","0110","0011","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0001","0001","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0101","0101","0111","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","0111","0111","0111","0110","0101","0101","0101","0100","0100","0111","0101","0100","0111","0111","0101","0110","0101","0111","0111","0111","0110","0110","0101","0100","0101","0110","0110","0101","0100","0100","0100","0110","0111","0111","0110","0011","0100","0111","0111","0111","0101","0100","0101","0111","0111","0110","0101","0101","0101","0100","0101","0110","0111","0111","0111","0111","0101","0011","0011","0101","0101","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0101","0110","0100","0011","0110","0111","0111","0111","0111","0111","0101","0101","0111","0111","0110","0110","0101","0101","0100","0100","0100","0101","0101","0100","0100","0100","0101","0101","0111","0111","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0100","0100","0111","0101","1001","1010","1010","0110","0110","1001","0011","1001","0110","0110","1001","0011","1001","0110","0110","1001","0100","1000","0101","0100","0100","0100","0101","0100","0101","0100","0011","0011","0100","0100","0011","0101","0110","0111","0110","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0101","0100","0100","0110","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0110","0101","0100","0100","0101","0100","0110","0110","0101","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0100","0101","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0110","0111","0110","0111","0111","0111","0110","0011","0011","0011","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","1000","1001","1001","1010","1011","1011","1100","1010","1001","1000","1000","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0101","0101","0110","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0010","0011","0011","0100","0100","0110","1000","1000","0110","0101","0101","0110","0111","1000","1000","1001","1000","1001","1011","1001","0111","1001","1000","1000","1000","0111","0110","0110","1000","1000","0111","0100","0011","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010"),
("0111","0111","0111","0111","0110","0110","0101","0011","0011","0010","0010","0011","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0010","0001","0001","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0111","0111","0100","0100","0110","0111","0110","0100","0101","0110","0111","0110","0100","0101","0110","0111","0110","0100","0110","0111","1000","0101","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0101","0101","0011","0101","0110","0101","0110","0101","0101","0101","0101","0101","0100","0100","0011","0011","0110","0011","0100","0110","0101","0101","0110","0111","0110","0100","0100","0100","0111","0111","0101","0100","0100","0101","0111","0110","0100","0101","0101","0101","0101","0101","0101","0110","0111","0111","0101","0011","0100","0100","0110","0110","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0101","0100","0011","0100","0101","0111","0111","0111","0111","0100","0011","0100","0110","0111","0111","0110","0110","0110","0101","0101","0101","0101","0100","0011","0011","0100","0011","0100","0101","0110","0110","0101","0110","0110","0110","0101","0101","1001","1011","1001","0110","0110","0101","0101","0101","0101","0110","1001","1010","1010","0110","0110","1001","0100","1001","0110","0110","1001","0100","1001","0110","0110","1001","0100","1000","0110","0110","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0110","0101","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0101","0101","0101","0100","0100","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0101","0101","0101","0101","0110","0111","0110","0110","0110","0111","0110","0110","0110","0110","0110","0111","0111","0111","0111","0110","0110","0100","0100","0101","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0010","0010","0010","0011","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0111","0111","0111","0111","0110","0011","0011","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","1000","1011","1001","1001","1011","1010","1010","1000","1000","0110","0110","0100","0101","0111","1010","1011","1011","1100","1100","1011","1001","1000","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0110","0110","0101","0011","0011","0110","0110","0101","0011","0101","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0100","0110","1000","1000","0110","0101","0110","0111","1000","1001","1001","1001","1000","1000","1010","1000","1001","1001","1001","1001","1000","1010","1001","1001","1000","0110","0110","0110","0111","1000","0111","0101","0100","0100","0011","0010","0010","0011","0100","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100"),
("0110","0101","0110","0101","0110","0111","0110","0101","0011","0010","0010","0010","0010","0011","0100","0011","0011","0011","0100","0011","0100","0100","0100","0011","0010","0011","0100","0011","0011","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0100","0101","0100","0100","0010","0100","0101","0101","0100","0010","0101","0101","0101","0100","0010","0101","0101","0101","0100","0011","0101","0101","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0011","0101","0110","0101","0110","0101","0100","0011","0011","0011","0011","0100","0011","0011","0101","0011","0101","0111","0101","0101","0110","0111","0110","0101","0100","0100","0110","0110","0101","0101","0100","0101","0111","0110","0100","0101","0110","0101","0101","0101","0101","0111","0111","0110","0100","0100","0101","0100","0101","0110","0010","0001","0001","0001","0001","0001","0001","0001","0011","0101","0100","0011","0100","0100","0101","0111","0111","0111","0101","0011","0100","0101","0110","0111","0111","0111","0110","0101","0101","0100","0101","0101","0011","0011","0011","0011","0011","0100","0101","0101","0110","0110","0110","0110","0110","0101","0110","1010","1011","1010","0111","0110","0101","0100","0100","0101","0101","1000","1011","1011","0111","0110","1010","0100","1010","0110","0110","1001","0100","0111","0101","0110","1001","0100","1000","0101","0100","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0100","0101","0101","0111","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0101","0101","0101","0101","0100","0101","0110","0110","0111","0111","0110","0111","0101","0100","0111","0111","0111","0111","0111","0110","0110","0110","0101","0101","0110","0101","0101","0110","0111","0110","0110","0110","0110","0110","0110","0101","0011","0100","0110","0110","0110","0110","0110","0110","0101","0100","0101","0101","0100","0100","0100","0100","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0101","0101","0101","0101","0011","0011","0011","0101","0101","0101","0101","0101","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","1000","1000","1001","0110","0110","0111","0111","0110","0101","1001","0100","0101","0011","0010","0011","1001","1010","1011","1011","1011","1100","1011","1001","1001","1010","1001","1010","1010","1010","1010","1001","1001","1001","1001","1001","1000","0110","0110","0100","0011","0100","0101","0110","0110","0110","0110","0111","0111","0110","0110","0110","0100","0011","0010","0011","0010","0010","0011","0010","0010","0010","0100","0101","0100","0111","1000","0111","0101","0110","0111","1001","0111","0100","0101","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0010","0010","0010","0100","0101","0011","0100","0101","0110","1000","1000","0110","0101","0101","0110","0111","1001","1000","0111","1001","1001","1000","0111","1000","1000","0111","1001","1000","0111","0111","1001","1010","1000","0111","1001","0111","0111","0110","0110","0111","1000","0111","0101","0100","0100","0011","0011","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0011","0100","0010","0010","0011","0011","0101","0011","0011","0011","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0110","0110"),
("0010","0010","0010","0011","0110","0111","0111","0111","0100","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0100","0010","0010","0001","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0001","0010","0010","0010","0010","0011","0010","0011","0011","0010","0100","0101","0011","0010","0011","0101","0101","0100","0010","0010","0110","0100","0011","0010","0011","0110","0011","0100","0011","0100","0110","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0101","0101","0100","0011","0011","0010","0010","0011","0100","0011","0011","0100","0100","0010","0100","0111","0101","0101","0110","0111","1000","0110","0100","0100","0110","0111","1000","0101","0100","0101","0110","1000","0110","0101","0111","0101","0101","0100","0101","0111","0111","0111","1000","0110","0101","0100","0101","0110","0010","0010","0010","0010","0001","0001","0010","0100","0101","0101","0110","0110","0101","0100","0101","0110","0111","0110","0110","0110","0101","0101","0110","0111","1000","0111","0110","0110","0101","0100","0100","0100","0011","0010","0010","0011","0100","0011","0100","0101","0110","0110","0100","0100","0101","0101","0100","0010","0011","0011","0101","0101","0011","0010","0010","0100","0110","1000","1001","1010","0111","0110","1001","0111","1001","1000","1000","1001","0011","0010","0101","1001","1010","1001","1001","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0101","0111","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0101","0101","0101","0100","0100","0101","0110","0111","0111","0111","0111","0110","0011","0010","0100","0111","0111","0110","0110","0110","0110","0110","0110","0101","0101","0110","0101","0111","0111","0111","0111","0110","0110","0110","0101","0011","0010","0011","0101","0111","0110","0110","0110","0101","0101","0100","0101","0101","0100","0101","0100","0101","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0101","0110","0111","1000","1000","1000","1000","1000","1000","1000","1000","1001","1010","0110","0100","0100","0010","0010","0110","0111","0111","0111","0011","0101","0010","0010","0011","0111","1000","1000","0111","0110","0101","0110","1010","1001","1001","1011","1010","1000","1000","1001","1001","1001","1001","1001","1001","1000","0110","0110","0100","0011","0100","0100","0101","0101","0101","0101","0101","0110","0110","0110","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0011","0100","0101","0111","0111","1000","0111","0111","1000","1000","1000","0111","0110","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0100","0100","0100","0011","0011","0011","0100","0011","0011","0100","0100","0100","0110","1000","1000","0110","0101","0101","0110","0111","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0101","0110","0111","1000","0111","0101","0011","0100","0100","0100","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0111","0111","1000","1000","0111","0111","0111","0111"),
("0010","0010","0100","0110","0110","0111","0111","0111","0101","0010","0010","0011","0100","0010","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0100","0110","0100","0011","0011","0110","0101","0101","0011","0011","0110","0100","0100","0011","0011","0110","0011","0100","0100","0100","0110","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0011","0100","0011","0011","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0101","0110","0101","0101","0110","0110","0111","0110","0100","0100","0101","0110","1000","0101","0100","0101","0110","0110","0110","0100","0110","0110","0101","0100","0101","0111","0111","0111","1000","0110","0100","0100","0101","0101","0010","0010","0010","0010","0010","0010","0011","0101","0100","0100","0101","0110","0101","0101","0101","0110","0110","0101","1000","1000","0101","0100","0101","0111","0111","0111","0111","0110","0110","0100","0100","0011","0010","0010","0001","0010","0010","0011","0100","0101","1000","1010","1001","0110","0011","0101","0111","0110","0110","0111","1001","0111","0011","0011","0100","0100","0101","0110","0101","0101","0101","0100","0101","0101","0100","0100","0101","0101","0011","0011","0011","0101","0101","0110","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0100","0011","0011","0110","0101","0101","0101","0100","0101","0110","0111","0111","0111","0111","0100","0011","0010","0001","0110","0111","0111","0110","0111","0111","0110","0110","0101","0101","0101","0110","0111","0111","0111","0111","0110","0110","0110","0100","0001","0010","0011","0100","0110","0110","0101","0110","0110","0101","0100","0101","0101","0101","0101","0101","0100","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0100","0111","0110","0110","0100","0011","0100","0101","0110","0110","0110","0110","0111","1001","1001","1001","1001","1010","1010","1010","1010","1010","1011","1010","0101","0011","0101","0010","0010","0111","1010","1001","0110","0101","0101","0100","0101","0101","0101","0100","0111","0100","0100","0010","0001","0100","1000","1010","1001","1010","1000","0100","0100","0101","0100","0100","0110","0011","0011","0100","0100","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0100","1000","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1001","0111","0101","0100","0110","0111","1000","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0111","0110","0101","0110","1000","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0111","1000","1000","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100"),
("0010","0011","0101","0101","0110","0111","0111","0111","0110","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0010","0001","0001","0010","0010","0001","0010","0010","0010","0011","0010","0001","0010","0010","0011","0011","0010","0100","0110","0101","0100","0011","0101","0110","0101","0100","0011","0101","0101","0100","0011","0011","0110","0100","0100","0100","0100","0110","0101","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0111","0101","0101","0110","0100","0110","0110","0100","0100","0101","0100","0111","0101","0100","0101","0100","0101","0110","0101","0101","0110","0110","0100","0101","0111","0111","0111","1000","0110","0100","0100","0101","0100","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0110","0101","0100","0101","0110","0110","0011","0111","1000","0101","0100","0101","0110","0111","0111","0111","0111","0110","0100","0100","0011","0011","0011","0001","0001","0010","0011","0011","0100","1000","1011","1010","1000","0101","1001","1010","1010","1010","1010","1010","1010","1000","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","0111","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0100","0100","0100","0100","0100","0011","0011","0010","0011","0011","0100","0100","0100","0100","0011","0100","0100","0011","0010","0010","0100","0110","0111","0101","0101","0101","0100","0101","0110","0111","0111","0111","0110","0100","0011","0001","0001","0011","0111","0111","0111","1000","0111","0111","0110","0110","0101","0101","0110","0111","0111","1000","1000","0111","0110","0110","0011","0001","0001","0011","0011","0101","0111","0110","0110","0101","0101","0100","0100","0100","0101","0110","0110","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0101","1000","0111","0100","0100","0100","0100","0101","0110","0101","0101","0111","1000","1001","1001","1000","0111","1010","1011","1011","1011","1001","1000","0111","0011","0110","0101","0100","0111","1001","1001","0110","0100","0101","0100","0100","0011","0101","0110","1001","0101","0101","0010","0010","0010","0010","0101","1010","1010","1011","1010","0110","0011","0101","0110","1001","0100","0100","0100","0101","0010","0001","0011","0101","0101","0100","0011","0011","0101","0110","0100","0011","0101","0111","0111","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1001","1001","1000","0111","0101","0111","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","0111","0111","0111","0111","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1001","1010","1001","1001","1000","1000","1000","1000","0111","1001","1010","1010","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","0111","0111","0111","0111","0111","0101","0110","0111","0111","0111","0110","0110","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101"),
("0011","0011","0011","0011","0100","0110","0111","0111","0101","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0101","0100","0101","0110","0100","0110","0110","0100","0100","0101","0100","0111","0101","0100","0101","0100","0101","0111","0101","0101","0110","0101","0101","0110","0111","0111","0111","0111","0101","0100","0100","0011","0010","0011","0010","0010","0010","0010","0101","0111","0110","0110","0110","0110","0111","0110","0100","0101","0110","0110","0100","0111","1000","0101","0100","0101","0110","0110","0111","0111","0110","0110","0101","0100","0011","0011","0010","0001","0010","0100","0110","0101","0101","1000","1011","1010","0111","1010","1101","1100","1011","1011","1101","1011","1100","1100","0111","0011","0100","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0011","0011","0011","0010","0010","0011","0011","0100","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0100","0100","0011","0011","0011","0100","1000","0111","0101","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0110","0110","0101","0100","0100","0100","0101","0110","0111","0111","0111","0110","0011","0011","0001","0001","0010","0110","0111","0111","1000","0111","0110","0110","0101","0101","0101","0101","0110","0110","0111","0111","0111","0110","0101","0001","0001","0001","0011","0100","0101","0111","0111","0110","0110","0100","0100","0100","0100","0100","0110","0101","0100","0100","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0001","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0101","1000","0100","0100","0100","0101","0101","0111","0111","0111","0111","1000","1001","1001","1000","1000","1000","1000","1010","1010","0111","0101","1000","0011","0100","0110","0100","0110","1001","1001","0111","0101","1000","0110","0101","0010","0011","0110","1001","0111","0110","0010","0101","0101","0100","0001","0101","1001","1010","1010","1100","0110","0100","0110","1001","0101","0100","0100","0101","0010","0010","0101","0011","0010","0110","0100","0101","0101","0011","0110","0100","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0110","0110","0110","0110","0111","0110","0110","0110","0111","0101","0110","0110","0101","0111","1000","0111","0111","0111","0111","0110","0101","0110","0101","0101","0101","0101","0101","0101","0110","0101","0110","0110","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100"),
("0011","0010","0011","0010","0100","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0110","0101","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0100","0110","0101","0101","0110","0101","0101","0101","0100","0100","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0100","0011","0100","0110","0111","0111","0110","0101","0101","0100","0010","0001","0010","0011","0011","0011","0010","0100","0110","0110","0110","0110","0101","0110","0101","0110","0101","0101","0110","0111","0100","0110","0111","0101","0100","0101","0110","0111","0111","0111","0110","0111","0101","0011","0010","0001","0001","0010","0011","0100","0100","0101","0110","0101","0110","1001","0111","1100","1100","1100","1011","1011","1101","1100","1011","1100","1011","0111","0110","0110","0111","0110","0110","1000","1000","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","1010","1001","1000","0110","0011","0011","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0110","0110","0100","0100","0100","0100","0101","0110","0110","0111","0111","0101","0100","0011","0010","0010","0010","0101","0111","0110","0111","0110","0101","0101","0101","0101","0101","0101","0110","0110","0110","0111","0110","0110","0101","0010","0010","0010","0010","0100","0101","0110","0110","0110","0101","0100","0100","0100","0100","0101","0110","0110","0100","0100","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0101","0011","0011","0100","0110","0111","1000","1000","1000","1000","1000","1000","1001","1001","0101","0110","0100","0101","0111","1000","0111","1001","0110","0110","0111","0101","1000","1001","1010","0111","0110","1001","0111","0101","0010","0010","0101","1001","0111","0101","0011","0100","0100","0010","0001","0011","0110","1010","1011","1000","1000","0111","0110","1001","0101","0100","0101","0101","0011","0010","0100","0001","0001","0101","0100","0110","0011","0001","0101","0101","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0100","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0111","0111","0110","0110","0110","0110","0101","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011"),
("0011","0010","0010","0010","0011","0101","0101","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0010","0001","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0101","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0111","0110","0100","0110","0110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0111","0101","0101","0110","0101","0110","0110","0100","0100","0101","0101","0111","0101","0100","0101","0101","0110","0110","0110","0110","0110","0110","0101","0110","0111","0111","0111","0111","0101","0011","0001","0010","0011","0011","0011","0011","0100","0110","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0111","0100","0110","0110","0100","0100","0101","0110","0110","0111","0111","0111","0111","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","1001","1011","1011","1100","1010","1011","1101","1100","1001","1100","1011","1000","0100","0011","0011","0011","0010","1001","1010","0100","0011","0100","0100","0100","0100","0101","0100","0100","0100","0100","0101","0100","0101","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0011","0011","0101","0111","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0010","0010","0011","0011","0011","0010","0011","0011","0011","0100","0011","0010","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0110","0111","0101","0100","0100","0100","0101","0110","0111","0111","0111","0101","0100","0011","0010","0010","0010","0100","0111","0111","0111","0110","0110","0101","0101","0101","0101","0101","0110","0110","0111","0111","0110","0110","0100","0001","0001","0001","0010","0100","0101","0110","0110","0110","0101","0100","0100","0101","0101","0101","0111","0110","0101","0101","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0101","1000","0111","0101","0100","0110","1001","0101","0010","0100","0100","0001","0101","0111","0111","0111","0111","1000","1001","1001","1001","1001","1001","0110","0101","1010","1000","0110","0010","0011","0110","1001","1000","0110","0101","0011","0101","0011","0001","0100","0110","0110","0101","1000","0011","0101","1000","1001","0101","0100","0100","0101","0010","0010","0010","0001","0001","0011","0100","0100","0010","0001","0011","0100","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0100","0100","0101","0101","0101","0101","0101","0100","0100","0110","0100","0101","0110","0101","0101","0110","0101","0101","0110","0100","0110","0110","0101","0110","0110","0101","0110","0101","0101","0110","0101","0101","0110","0101","0101","0110","0101","0110","0110","0101","0110","0110","0101","0110","0110","0101","0110","0110","0101","0110","0110","0110","0111","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0100","0100","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0010","0011","0010","0100","0101","0011","0011","0010","0100","0110","0100","0011"),
("0111","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0010","0010","0001","0010","0100","0011","0010","0010","0010","0010","0011","0011","0010","0001","0001","0010","0010","0010","0010","0011","0100","0011","0011","0110","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0101","0101","0010","0100","0101","0110","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0011","0100","0111","0101","0101","0110","0101","0110","0110","0100","0100","0101","0100","0111","0101","0100","0101","0101","0110","0110","0111","1000","0111","0111","0111","0110","0110","1001","1001","0110","0101","0100","0011","0011","0100","0011","0011","0011","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0110","0110","0111","0100","1000","0111","0101","0100","0101","0110","0110","0111","0111","0110","0100","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0101","1010","1011","1011","1011","1001","1011","1100","1100","1001","1010","1011","1010","0101","0010","0010","0010","0010","0110","0110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0011","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","1000","0111","0110","0111","0111","0110","0111","0111","0111","0110","0100","0010","0010","0010","0001","0001","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0101","0100","0100","0111","0111","0101","0100","0100","0100","0101","0110","0111","0111","0111","0101","0100","0011","0010","0010","0010","0100","0111","1000","1000","0111","0110","0110","0101","0101","0101","0101","0110","0111","0111","0111","0111","0110","0100","0001","0001","0001","0010","0100","0101","0110","0110","0110","0101","0100","0100","0101","0101","0101","0111","0110","0100","0101","0011","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0101","0110","0101","0101","0110","0101","0101","0101","0100","1000","1000","0101","0010","0010","0110","0010","0101","0111","0101","0101","0101","0101","1000","1000","0111","0110","0101","0101","0101","1010","1000","0111","0010","0011","0111","1001","1001","0110","0100","0001","0110","0011","0001","0100","0110","0100","0010","0101","1001","0100","1001","1010","0101","0100","0100","0101","0010","0010","0010","0001","0001","0011","0100","0100","0010","0001","0010","0100","0101","0110","0110","0101","0101","0101","0110","0110","0101","0101","0101","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0110","0111","0110","0110","0101","0101","0101","0110","0101","0101","0101","0101","0110","0101","0100","0110","0111","0100","0100","0111","0100","0100","0110","0110","0110","0110","0101","0011","0100","0110","0011","0011","0101","0110","0110","0100","0011","0101","0101","0011","0100","0110","0110","0101","0011","0011","0101","0100","0011","0101","0101","0101","0100","0011","0100","0101","0011","0100","0101","0101","0101","0100","0100","0100","0100","0011","0100","0101","0101","0100","0100","0101","0100","0100","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0101","0011","0011","0010","0100","0110","0100","0011","0011","0100","0110","0110","0011","0100","0011","0110","0111","0100","0101","0011","0110","0111","0101","0100"),
("1001","0111","0100","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0100","0101","0100","0011","0011","0011","0011","0011","0001","0010","0100","0100","0011","0010","0010","0011","0100","0100","0010","0001","0010","0100","0011","0010","0001","0011","0100","0011","0010","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0100","0110","0011","0010","0011","0110","0110","0110","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0100","0100","0111","0101","0101","0110","0101","0110","0110","0011","0100","0110","0101","0111","0101","0100","0101","0101","0101","0111","0111","0111","0110","0110","0111","1001","0111","0110","0110","0100","0101","0110","0110","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0101","0110","0110","0101","0101","0101","0101","0101","0110","0100","1000","0111","0100","0100","0101","0110","0110","0111","0110","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0110","1010","1010","1010","1011","1000","1010","1011","1011","1001","1010","1010","1010","1000","0011","0010","0010","0010","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0110","0110","0110","0100","0011","0011","0011","0100","0100","0101","0100","0101","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0100","0101","0101","0100","0111","1000","0110","0100","0100","0100","0110","0110","0111","0111","0111","0110","0100","0011","0001","0001","0010","0100","0111","1000","1000","0111","0110","0110","0101","0101","0101","0110","0111","1000","0111","0111","0111","0110","0011","0001","0001","0001","0010","0100","0101","0110","0110","0101","0101","0101","0100","0101","0101","0101","0111","0110","0100","0101","0011","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0111","1001","1001","1000","0101","0100","0111","1001","1001","1001","1000","0100","0011","0110","0111","0111","1001","1000","1010","1010","1001","1010","1011","1010","1010","1001","0111","0101","1010","0111","0111","0010","0011","0111","1001","1001","0111","0011","0001","0101","0011","0001","0100","0111","0011","0011","0011","0111","1010","1000","1011","0110","0100","0100","0101","0010","0010","0010","0001","0001","0011","0100","0100","0010","0001","0010","0100","0100","0111","0111","0101","0011","0011","0110","0111","0100","0011","0100","0111","0111","1000","0110","0101","0010","0010","0011","0011","0101","0111","1000","0111","0110","0100","0010","0011","0111","0110","0011","0010","0101","0101","0110","0100","1000","1001","0100","0010","1000","0011","0010","1000","1001","1001","1001","0110","0001","0011","0111","0010","0010","0111","1000","1000","0011","0001","0110","0101","0001","0100","1000","1000","0110","0001","0010","0111","0011","0010","0110","1000","1000","0011","0001","0101","0110","0001","0010","0111","1000","0111","0010","0010","0110","0101","0001","0011","0111","0111","0111","0111","0110","0010","0101","0110","0010","0100","1000","0111","0111","0110","0011","0100","0011","0101","0111","0101","0100","0011","0101","1000","0100","0101","0011","0110","0111","0110","0100","0100","0101","0111","0111","0100","0101","0100","0111","1000","0101","0101","0100","0110","1000","0110","0101"),
("0100","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0011","0010","0010","0100","0101","0100","0010","0010","0011","0100","0011","0010","0001","0011","0101","0011","0011","0010","0011","0011","0011","0001","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0101","0011","0011","0011","0110","1000","0111","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0101","0011","0101","0110","1001","1001","0110","0101","0110","0110","0011","0110","1100","1000","0111","0101","0100","0111","1001","0101","0111","1011","0111","0100","0100","0101","0111","0101","0011","0011","0011","0011","0110","1001","0111","0111","1000","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0100","1000","0111","0100","0100","0101","0110","0110","0110","0110","0101","0011","0011","0010","0001","0010","0010","0010","0010","0100","0101","0010","0010","0011","0101","0110","1001","1010","1010","1011","0111","1001","1011","1011","1000","1000","1010","1010","1000","0011","0010","0010","0010","0110","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","1000","0111","0111","0111","0111","0111","0110","0111","0110","0111","0110","0110","0111","0111","0111","0111","0101","0101","0101","0110","0100","0011","0011","0011","0110","0111","0111","0111","0111","1000","0111","0111","0100","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0101","0101","0011","0110","1000","0110","0101","0101","0101","0101","0110","0111","0111","0111","0110","0100","0011","0001","0001","0010","0100","0111","1000","1000","0111","0110","0110","0101","0101","0110","0110","0111","0111","0111","0111","0111","0110","0100","0001","0001","0001","0010","0100","0100","0110","0110","0101","0101","0101","0100","0100","0101","0101","0111","0110","0100","0101","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0100","0101","0100","0101","0011","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0111","0111","0110","0101","0101","1000","0111","0111","1001","0111","0100","0011","0011","0111","1001","1010","1010","1011","1011","1011","1011","1100","1011","1011","1010","0110","0101","1010","1000","0111","0011","0011","0111","1001","1000","0111","0011","0001","0110","0011","0001","0101","0111","0101","0011","0101","0101","1001","1010","1010","1011","0101","0100","0101","0010","0010","0010","0010","0001","0011","0100","0100","0010","0001","0010","0100","0101","1001","1000","0110","0011","0011","0110","0111","0100","0011","0100","0111","0110","0101","0110","0101","0011","0011","0011","0011","0101","0110","0110","0111","0111","0100","0010","0100","0111","0110","0011","0011","0101","0111","1000","0101","1000","1001","0100","0010","1000","0100","0010","1000","1001","1001","1001","0110","0010","0100","1000","0010","0010","0111","1001","1001","0011","0010","0110","0110","0010","0100","1001","1001","0111","0010","0011","1000","0100","0010","0110","1001","1001","0100","0010","0101","0111","0010","0011","1000","1001","1000","0011","0010","0111","0101","0010","0100","1000","1000","1000","1000","0111","0001","0100","0111","0001","0101","1000","1000","1000","0110","0100","0101","0100","0101","1000","0110","0101","0100","0101","1000","0101","0101","0100","0111","1000","0111","0101","0100","0101","1000","1000","0100","0110","0100","0111","1000","0101","0101","0100","0111","1000","0110","0101"),
("1010","1010","1010","1010","1000","0100","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0101","0100","0011","0100","0101","0110","0100","0011","0011","0100","0100","0100","0011","0011","0100","0110","0100","0011","0011","0100","0100","0100","0011","1000","0110","0010","0010","0010","0010","0011","0011","0011","0011","0100","0011","0101","0110","0100","0101","0101","0110","1000","1001","1010","1010","1001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0110","1011","1000","0011","0110","0011","0011","0101","1001","1010","0110","0101","0110","0110","0101","0111","1001","0111","0111","0101","0111","1001","1010","1000","0110","1010","0110","0011","0011","0011","0011","0011","0011","0100","0100","0011","0111","1011","1010","1010","1011","0111","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","1000","0111","0100","0100","0101","0101","0110","0110","0110","0101","0100","0101","0011","0011","0100","0100","0011","0011","0100","0100","0100","0100","0101","0101","0110","1001","1001","1001","1010","0110","1000","1010","1010","1000","1000","1001","1001","1000","0100","0010","0010","0010","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0111","0111","0111","1000","1000","1000","0111","0111","0101","0011","0011","0100","0110","0111","1000","1000","0101","0011","0011","0011","0010","0100","0101","0101","0101","0101","0101","0110","0110","0110","0111","0111","0011","0100","0100","0101","0100","0011","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0100","0100","0100","0100","0101","0101","0011","0110","0111","0101","0100","0101","0101","0101","0110","0111","0111","0111","0110","0101","0011","0001","0010","0010","0100","0111","1000","1000","0111","0111","0110","0101","0101","0110","0110","0111","0111","0111","0111","0111","0110","0011","0001","0001","0001","0011","0101","0101","0110","0110","0101","0110","0101","0101","0101","0101","0101","0111","0110","0100","0101","0100","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0001","0100","0100","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0101","0101","0110","1001","0111","1010","0111","0101","0100","0100","0100","0100","1000","1000","1000","1010","1011","1011","1011","1011","1011","1011","1010","0110","0111","1010","1001","1000","0110","0110","0110","1010","0111","0110","0011","0100","0110","0100","0100","0111","1000","0110","0011","0100","0011","0100","1001","1010","1000","1010","0100","0101","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0101","1001","1001","0110","0011","0100","0110","1000","0100","0100","0100","0110","0110","0101","0101","0110","0011","0011","0011","0011","0101","0101","0101","0101","0111","0101","0011","0100","0111","0110","0011","0011","0101","0111","1000","0101","1001","1010","0100","0001","1000","0100","0010","1001","1010","1010","1001","0111","0010","0100","1000","0011","0011","1000","1001","1001","0011","0011","0110","0110","0010","0100","1001","1001","0111","0010","0011","1000","0100","0010","0111","1001","1001","0101","0100","0110","0111","0011","0100","1001","1001","1001","0011","0100","0111","0110","0011","0101","1001","1001","1001","1000","0111","0001","0100","0111","0001","0100","1001","1001","1000","0110","0100","0101","0100","0111","1000","0111","0100","0100","0110","1000","0101","0110","0101","0111","1000","0111","0101","0101","0101","0111","1000","0100","0110","0100","0111","0111","0101","0101","0100","0101","0101","0101","0101"),
("1100","1011","1011","1011","1011","1001","0100","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0011","0110","1001","1001","1001","1001","1001","1000","1010","1001","1010","1010","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0111","1001","1001","0111","1000","1000","1001","1001","1010","1010","1010","1011","1000","1010","1001","1000","0111","1000","0111","0110","1000","1001","1001","0111","0010","0011","0100","0011","0011","0100","0100","0101","0101","0101","0110","0110","1000","1100","1011","1001","1100","1001","1000","1001","1000","1000","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1010","1010","1001","1001","1000","0101","0011","0011","0110","0110","0110","0111","0111","0111","0111","0111","1001","1010","1001","1010","1010","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0100","0100","0011","0011","0101","0101","0101","0110","0100","0101","0110","0110","0101","0110","0101","0101","0101","0011","0010","0010","0010","0100","0100","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0101","0110","0110","0110","0110","0101","0101","0100","0011","0010","0010","0010","0011","0011","0101","0111","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0010","0001","0100","0111","0110","0100","0111","1000","1001","1000","0100","0011","0011","0010","0010","0100","0110","0101","1001","1000","0111","0111","0111","0111","0101","0010","0011","0101","0100","0100","0111","1010","1000","0101","0100","0010","0110","1000","0110","0101","0101","0101","0101","0110","0111","0111","0111","0110","0101","0100","0001","0010","0010","0100","0111","1000","1000","0111","0111","0110","0101","0101","0110","0110","0111","1000","1000","0111","0111","0110","0100","0001","0001","0001","0011","0100","0100","0110","0110","0110","0101","0101","0110","0101","0101","0110","1000","1001","0110","0100","0100","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0100","0101","0100","0100","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0001","0010","0010","0001","0011","0111","1001","1010","1001","1010","1010","0111","0101","0110","0111","0111","0111","1000","1010","1001","1011","1011","1011","1011","1011","1011","1010","1000","0101","0111","1010","1000","0111","0110","0111","1000","1010","1001","0111","0110","0110","1000","0101","0111","0111","0111","1000","0101","0101","0101","0101","0110","1011","0111","1001","1000","0100","0010","0011","0011","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","1000","0111","0110","0011","0100","0110","1000","0101","0100","0101","0111","1000","1000","0110","0110","0011","0011","0100","0100","0101","0111","1000","0110","0111","0101","0011","0100","0111","0111","0011","0100","0101","0110","1000","0101","1000","1010","0100","0010","1000","0100","0010","1000","1001","1001","1001","0110","0010","0100","1000","0011","0011","0111","1001","1001","0011","0010","0111","0110","0010","0100","1001","1001","0111","0010","0011","1000","0100","0010","0111","1001","1001","0100","0100","0110","0111","0011","0100","1001","1001","1001","0011","0100","0111","0110","0100","0101","1001","1001","1001","1001","1000","0001","0100","0111","0001","0100","1001","1001","1001","0111","0100","0101","0101","0110","1000","0110","0100","0100","0100","0111","0101","0110","0110","0111","0111","0111","0101","0110","0110","0111","0110","0011","0011","0011","0110","0110","0101","0100","0001","0000","0001","0010","0100"),
("1010","1010","1001","1001","1001","1001","0111","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0100","0110","1000","1000","1001","1001","1001","1010","1000","0100","0010","0010","0011","0101","0100","0010","0101","1010","1010","1010","1000","0110","1000","1010","0111","0110","1010","1010","1010","1010","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","0111","0101","0110","1001","1011","1010","1010","1001","1001","1001","1001","1000","0111","1000","1001","1000","1001","1000","1000","0110","0101","0100","0011","0010","0010","0011","0011","0101","1000","0111","0101","1000","1010","1010","1010","0111","0110","1000","1000","0110","0110","0111","1000","1010","1010","1001","1010","1001","1010","1011","1010","1010","1010","1010","1010","1011","1100","1011","1010","1010","1010","1001","0111","0101","0111","1001","1001","0110","0110","0110","1000","1000","1010","1000","0100","0101","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0011","0110","1000","1000","1000","1000","0100","0111","1001","1000","0110","0101","1000","0111","0111","0100","0010","0010","0010","0101","0111","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0100","0101","0101","0110","0110","0110","0111","0110","0101","1000","0111","1000","1000","0111","1000","1010","1010","1010","1000","0110","0101","0010","0010","0100","0101","0101","0101","0100","0100","0100","0101","0100","0011","0101","0011","0010","0100","0101","0100","1000","1000","0111","0110","0101","0110","0100","0011","0011","0011","0010","0001","0010","0110","0111","0110","0011","0100","1000","1001","0110","0101","0101","0101","0101","0110","0111","0111","0111","0110","0101","0011","0001","0010","0010","0011","0111","1010","1010","1001","1000","0111","0111","0110","0111","0111","1000","1000","1001","1001","1001","0111","0100","0001","0001","0001","0010","0100","0100","0110","0110","0101","0101","0100","0011","0100","0011","0100","0101","0101","0101","0100","0100","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0001","0010","0011","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0011","0111","0111","0110","0100","0101","0111","0100","1000","1001","1001","1001","1001","1011","1010","1011","1011","1010","1010","1010","1011","1011","0111","0100","0100","0111","0110","0111","0101","0101","0110","0111","0111","0111","0110","0110","0101","0111","0111","0111","0101","0101","0101","0101","0101","0101","0101","1000","1011","1010","1011","1000","0011","0011","0100","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","1000","0111","0110","0100","0101","0111","1000","0101","0100","0110","0111","0111","1000","0110","0110","0100","0100","0100","0100","0101","0111","0111","0111","0111","0101","0011","0100","1000","0111","0100","0100","0101","0110","0111","0101","1000","1001","0111","0111","1000","0111","0111","1000","1001","1001","1001","1000","0111","0111","1001","0110","0110","1000","1001","1001","0110","0110","1000","0111","0110","0110","1001","1001","0111","0101","0110","1000","0101","0100","0111","1001","1001","0110","0110","0111","1000","0110","0110","1001","1001","1000","0101","0101","1000","0110","0101","0110","1001","1001","1000","1000","1000","0100","0101","0111","0100","0101","1000","1000","1000","0111","0101","0110","0101","0101","0111","0111","0011","0001","0001","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0001","0010","0101","0101","0100","0011","0001","0000","0001","0010","0101"),
("0110","0111","0111","0110","0110","0110","0110","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","1000","1010","1010","1010","1010","1010","1010","1001","0101","0011","0100","0101","0100","0100","0100","0101","0101","0110","0100","0010","0011","0011","0010","0010","0100","0110","0110","0101","0101","0101","0110","0110","0110","0110","0101","0110","1011","1101","1100","1101","1100","1011","1100","1001","0100","0101","0101","0100","0100","0101","0101","0101","0101","1001","1011","0101","0100","1000","1010","0111","0011","0010","0010","0010","0011","0100","0101","0011","0010","0100","0111","0110","0110","0011","0011","1000","1011","1010","1001","1001","1010","1001","0101","0100","0100","0100","0110","1010","1011","1010","1001","0111","1000","1001","1100","1010","1001","1001","1001","0111","0110","0101","0101","0110","0110","0100","0101","0011","0100","0110","0110","0101","0100","0011","0010","0100","0100","0100","0100","0100","0011","0100","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","1010","1000","0100","0100","0110","0101","1001","1011","1011","1011","1100","0111","1010","1100","1100","1010","1000","1011","1010","1001","0110","0011","0010","0011","0100","0110","0110","0011","0010","0010","0010","0111","1001","1001","1001","1000","1001","1000","1000","0111","0110","1001","1010","1010","1010","1010","1010","1010","1010","1000","0110","1000","1000","0111","0101","1000","1000","1000","0111","0101","0011","0011","0011","0010","0010","0011","0011","0011","0100","0100","0011","0010","0011","0011","0011","0100","0011","0100","0110","0101","0011","0011","0011","0011","0010","0010","0100","0011","0100","0100","0011","0011","0010","0010","0100","0101","0100","0010","0010","0100","0100","0011","0011","0011","0011","0100","0110","0110","0111","0111","0110","0101","0011","0010","0010","0010","0100","0111","0110","0110","0101","0100","0100","0011","0011","0100","0011","0100","0100","0101","0101","0100","0101","0100","0010","0010","0010","0010","0100","0100","0110","0110","0110","0101","0100","0011","0011","0011","0100","0100","0100","0100","0100","0101","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0011","0011","0011","0110","0011","0111","1000","1001","1010","1010","1010","1001","1010","1011","1011","1011","1010","1010","1010","1011","1010","1000","0011","0011","1000","0110","0111","0101","0100","0111","0110","0110","0110","0110","0111","0111","1000","0111","0111","0101","0101","0101","0101","0100","0100","0100","0101","0111","0111","0100","0101","0011","0010","0100","0100","0101","0101","0101","0101","0101","0101","0110","0101","0100","0101","0100","0011","0100","0100","0101","0101","0100","0100","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0110","0101","0100","0101","0110","0110","0100","0100","0100","0101","0111","0100","0110","0111","0111","0111","0110","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","0111","1000","1000","0110","0111","1000","1000","0111","0111","1000","1000","0111","0111","0111","0111","1000","1000","0111","0111","0111","0110","0110","0010","0011","0011","0001","0000","0000","0001","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0000","0000","0001","0011","0100","0011","0100","0001","0000","0000","0010","0100"),
("0111","0111","0111","0111","0111","0111","1000","0110","0001","0010","0100","0101","0101","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0100","0100","0100","0101","0111","1001","1001","1001","1001","1001","1001","1001","0110","0101","0101","0101","0101","1000","1001","1001","1000","0110","0011","0010","0011","0010","0001","0011","1001","1001","0100","0100","0011","1000","1001","1001","1001","1000","1000","1010","1010","1010","1010","1010","1001","1001","1001","0101","0111","1000","0100","0100","0101","0100","0100","0100","1001","1011","0100","0011","1001","1011","1001","0100","0011","0011","0100","0100","0011","0100","0100","0100","0100","0011","0011","0100","0101","0111","1011","1100","1100","1100","1100","1011","1011","1000","0011","0010","0100","0101","0100","0110","1000","1001","1000","1001","1001","1011","1011","0110","0101","0111","0100","0001","0001","0010","0011","0101","0101","0101","0101","0101","0011","0001","0100","0101","0101","0101","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0101","0100","0100","0100","0011","0101","0111","0111","1010","1100","1100","1011","1100","1001","1011","1101","1100","1011","1001","1011","1011","1010","1000","0101","0100","0100","0011","0110","0110","0110","0100","0100","0100","0111","1000","0111","1000","1000","1000","1001","1001","1000","0111","1001","1001","1001","1001","1000","1000","1000","1000","0111","0110","0111","0110","0011","0010","0110","0110","0100","0011","0010","0011","0011","0100","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0100","0011","0011","0011","0100","0011","0011","0011","0010","0101","0110","0111","0111","0111","0110","0101","0101","0110","0110","0101","0101","0100","0001","0010","0100","0110","0101","0100","0100","0011","0100","0110","0110","0110","0111","0110","0101","0100","0001","0010","0010","0100","0111","0101","0101","0100","0100","0100","0011","0011","0100","0011","0100","0101","0101","0101","0100","0101","0100","0001","0001","0001","0010","0100","0101","0110","0110","0110","0101","0100","0100","0100","0100","0101","0110","0101","0100","0100","0101","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0010","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","1000","1000","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1010","1011","1010","1000","0011","0011","0111","0110","1000","0111","0110","1001","1000","1001","1001","1001","1010","1010","1001","1000","1000","0111","0100","0100","0100","0101","0101","0110","0100","0011","1000","0010","0010","0011","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0011","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0101","0110","0110","0101","0101","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0010","0010","0011","0001","0000","0000","0010","0011","0011","0010","0011","0011","0011","0100","0011","0011","0011","0011","0000","0000","0000","0010","0011","0010","0011","0001","0001","0001","0001","0001"),
("1011","1010","1010","1010","1010","1010","1001","1010","0111","0011","0101","0101","0100","0101","0110","0101","0101","0101","0110","0110","0101","0110","0111","0101","0110","0101","0110","0110","0110","0110","0011","0100","0101","0101","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0101","0100","0101","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","0011","0100","0110","0101","0100","0101","1010","1010","0100","0101","0100","1001","1011","1010","1010","1010","0110","0100","0110","0111","0111","0111","1000","1000","1001","1000","1010","1010","0110","0111","1000","0111","0110","0110","0110","1000","0100","0011","1010","1100","1001","0100","0100","0100","0101","0100","0100","0011","0100","0100","0100","0011","0011","0011","0101","0111","0111","1000","0111","0111","0111","1000","1000","1000","0100","0010","0100","0101","0100","0011","0110","1010","1010","1010","1010","1011","1000","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0100","0011","0011","0010","0011","0101","0110","0111","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0101","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0101","0100","0100","1000","0111","0111","1010","0110","0101","0110","1001","1010","1011","1011","1011","1100","1000","1010","1100","1100","1011","1000","1001","1011","1010","1001","1000","1000","0110","0101","1010","1000","1010","1000","1000","1000","0111","0111","0111","0101","0010","0011","0111","1000","0111","0110","1000","1000","1000","1000","1000","1000","1000","1000","0111","0011","0011","0010","0001","0010","0011","0011","0011","0011","0010","0011","0011","0010","0011","0101","0101","0101","0011","0010","0100","0110","0100","0011","0010","0010","0011","0011","0010","0011","0101","0100","0100","0011","0001","0010","0011","0100","0111","0101","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0110","0111","0101","0101","0101","0100","0101","0110","0111","0111","0111","0110","0101","0100","0001","0010","0010","0100","0111","0111","0111","0110","0101","0101","0100","0100","0101","0100","0101","0101","0110","0111","0110","0110","0100","0001","0001","0010","0010","0100","0101","0111","0110","0110","0101","0100","0100","0100","0101","0101","0110","0101","0100","0100","0101","0011","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0010","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0101","1000","1001","1011","1010","1010","1001","1010","1001","1001","1011","1010","1011","1000","0100","0110","1001","1010","1010","1010","1011","1011","1011","1010","1000","1011","1011","1011","1100","1011","1011","1011","1000","0100","0111","1000","0101","0101","0101","0101","0111","0110","0010","0001","0111","0110","0001","0110","0010","0011","0100","0100","0100","0011","0100","0101","0110","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0111","1001","1010","1001","1010","1010","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0100","0110","1000","1000","0111","0111","1000","1000","1000","1000","0111","1000","1000","0101","0101","0101","0111","1000","0111","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0010","0010","0010","0010","0010"),
("0100","0100","0100","0011","0100","0011","0011","0011","0011","0010","0100","0100","0010","0101","0110","0010","0010","0011","0110","0100","0011","0101","0101","0011","0100","0100","0011","0010","0010","0100","0011","0100","0011","0011","0011","0011","0100","0100","0011","0011","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0011","0011","0101","1000","1001","1001","1001","1001","0111","0111","0101","1010","1011","1011","1011","1011","0110","0001","0010","1000","1011","1100","1011","1011","1011","1100","1011","1000","0101","0101","0100","0101","0101","0101","0101","0101","0110","0111","1010","1011","1001","0100","0011","0100","0100","0100","0100","0010","0011","0100","0100","0011","0010","0001","0111","1000","0011","0100","1000","1010","1010","1010","1010","1011","1001","0101","0100","0101","0101","0100","0101","0101","0101","0110","0110","0110","0101","0101","0101","0101","0100","0100","0100","0011","0001","0010","0100","0100","0101","0110","0111","0110","0101","0100","0100","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0101","0100","0110","1011","1010","1010","1011","0110","0011","0100","1001","1010","1001","1010","1010","1001","0100","0111","1001","1001","1001","0101","0100","1000","1000","1000","1000","0110","0110","0111","1011","1011","1011","1000","0101","0101","1000","1001","1000","0101","0010","0011","0110","0111","0110","0101","1000","1001","1001","1001","1000","1000","1000","1000","0110","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0100","0111","1000","0110","0110","0100","0100","0100","0110","1000","0110","0100","0101","0110","0111","0110","0110","0111","0110","0111","0111","0110","0100","0011","0011","0100","0111","0100","0010","0010","0010","0010","0011","0010","0010","0001","0010","0110","1000","0110","0101","0101","0100","0101","0110","0111","0111","0111","0110","0101","0100","0001","0010","0010","0100","0111","0111","1000","0110","0110","0110","0101","0101","0110","0101","0110","0110","0111","0111","0111","0110","0100","0001","0001","0001","0010","0100","0101","0110","0110","0110","0101","0100","0100","0100","0100","0101","0110","0110","0100","0100","0100","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0100","0100","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0111","1001","1001","1010","1000","0110","0100","0101","0101","1000","0110","0111","0001","0010","0110","1010","1011","1011","1011","1100","1011","0110","0110","1001","1001","1001","1000","1001","1010","1000","0111","0100","0101","0111","0011","0011","0100","0110","0111","0111","0101","0011","0101","1010","0100","1000","0101","0100","0010","0001","0101","0100","0110","0100","0001","0110","0101","0100","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0110","0110","0110","0110","0110","0101","0110","0101","0101","0110","0100","1000","1010","1010","1010","1010","1010","1001","1001","1001","0111","0111","0111","1000","1000","1000","1000","0111","0111","0111","0111","0011","0011","0011","0011","0011","0100","0110","0110","0110","0011","0011","0011","0011","0011","0101","0110","0110","0101","0011","0011","0011","0011","0011","0110","0110","0111","0111","0111","0111","0110","0101","0110","0111","0111","0111","1000","1001","1000","1001","1001","1000","1000","1000","0110","0101","0101","0110","1000","0100","0010","0010","0010","0010","0010","0001","0010","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0100","0110","0101"),
("0001","0001","0011","0010","0011","0010","0010","0010","0001","0001","0100","0101","0100","0100","0100","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0011","0100","0011","0011","0100","0100","0101","0100","0011","0011","0100","0011","0011","0011","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0101","0100","0100","0110","0110","1001","1001","1001","1001","1001","1010","1001","1001","1001","1000","0111","0101","0001","0010","0010","0011","0101","0101","0110","0110","0101","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0100","0110","1011","1100","1100","1011","1001","1001","1001","1000","1000","1000","0111","0111","1000","0111","0111","0110","0111","1000","0011","0001","0001","0110","1011","1011","1010","1010","1010","1001","0111","0101","0101","0110","0100","0011","0011","0011","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0010","0100","1000","1000","1000","1000","0111","1000","0101","0100","0100","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0011","0011","0100","0101","0101","0110","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0110","0111","0110","0101","1000","1011","1100","1000","0100","0111","1001","0101","0100","0110","1010","1011","0101","1000","0111","0100","0101","0111","0101","1011","1011","0111","0100","0101","1000","1000","1010","1010","1001","0011","0001","0100","0101","0100","0100","0011","0010","0010","0010","0011","0010","0010","0110","0110","0110","0101","0100","0101","0101","0100","0100","0011","0100","0011","0011","0100","0100","0011","0011","0011","0011","0101","0101","0101","0111","0111","0111","1000","1001","1001","1001","1001","1000","0111","0111","0111","0111","0110","0110","0110","0111","0110","0101","0101","0101","0101","0100","0011","0010","0101","0111","0010","0010","0010","0010","0010","0010","0001","0010","0001","0110","1000","0110","0101","0101","0100","0101","0110","0111","0111","0111","0110","0100","0100","0001","0001","0010","0100","0111","0111","1000","0110","0110","0110","0101","0101","0110","0101","0101","0110","1000","1000","0111","0110","0100","0001","0001","0001","0010","0101","0101","0110","0101","0101","0101","0101","0100","0100","0101","0101","0110","0110","0100","0100","0100","0100","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0110","0111","1001","1000","1011","0110","0100","0100","0011","0111","0110","1000","0100","0010","0111","1010","1011","1010","1011","1010","1001","0100","0101","0101","0101","0010","0010","0101","0100","0101","0011","0101","0100","0100","0011","0100","0110","0111","0101","0010","0100","0011","0100","1001","1000","1001","1000","0101","0011","0001","0101","0100","0110","0011","0001","0100","0101","0100","0110","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0100","1000","1010","1010","0111","0110","0110","1001","1010","1010","1000","1000","1000","0110","0110","0110","0110","0111","1000","1000","1000","0100","0100","0100","0100","0100","0101","0101","0110","0100","0011","0100","0100","0011","0100","0100","0101","0101","0011","0100","0100","0011","0011","0100","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1001","1000","1000","1000","0111","1000","1001","0110","0110","0111","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0101","1000","0110"),
("0010","0011","0011","0011","0011","0011","0011","0010","0001","0001","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0101","0011","0011","0010","0010","0001","0001","0010","0010","0011","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0101","0101","0101","0011","0101","0101","0100","0100","0100","0110","0101","0101","0110","0101","0110","0010","0010","0011","0101","0100","0011","0010","0011","0011","0011","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1001","1001","1001","1001","1010","1010","1101","1101","1101","1100","1100","1100","1100","1101","1101","1101","1001","0010","0001","0010","0011","0010","0011","0011","0011","0011","0011","0011","1000","1101","1101","1101","1010","0111","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0110","0110","0100","0010","0100","1001","1001","1000","1000","1000","0111","0101","0011","0100","0101","0110","0110","0110","0110","0110","0110","0100","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0100","0011","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0110","0001","0000","0010","0111","1001","1000","0111","0111","0011","0010","0010","0010","0101","1001","0101","1000","0011","0010","0001","0100","0101","1000","0111","0011","0010","0010","0101","0101","0101","0101","0011","0010","0001","0010","0010","0010","0011","0011","0011","0011","0011","0100","0100","0101","0110","0110","0111","0111","1000","1001","1010","1011","1011","1001","1001","0111","0011","0100","0101","0011","0011","0011","0100","0100","0011","0100","0011","0011","0010","0011","0100","0100","0101","0100","0100","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0110","1000","0110","0101","0101","0101","0101","0110","0111","0111","0111","0110","0100","0100","0001","0010","0010","0100","0111","1000","1000","0110","0110","0110","0101","0101","0110","0101","0110","0111","0111","0111","0111","0111","0100","0001","0001","0001","0010","0101","0101","0110","0110","0110","0110","0101","0100","0100","0101","0101","0110","0110","0100","0100","0100","0100","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0111","0111","1001","1001","0110","0100","0110","0111","1000","1000","1000","0011","0111","0111","0111","0110","1000","0110","0111","0011","0110","0101","0101","0001","0011","0111","0110","0100","0010","0010","0101","0011","0110","0111","0110","0100","0010","0010","0010","0011","0011","0110","1010","0111","1001","0110","0011","0001","0101","0100","0111","0100","0001","0101","0110","0100","0101","0101","0101","0100","0010","0010","0010","0011","0011","0101","0101","0101","0101","0101","0100","0010","0011","0011","0010","0100","0101","0101","0101","0100","0101","0100","0010","0010","0010","0010","0100","0101","0101","0101","0101","1000","1001","1010","0101","0010","0010","1000","1010","1001","1001","1001","1001","0110","0110","0010","0101","0111","1001","1001","1000","0101","0110","0011","0010","0010","0101","0110","0110","0100","0101","0101","0010","0001","0010","0110","0110","0101","0100","0101","0100","0001","0001","0100","0111","1000","1000","0110","0100","0100","0101","0100","0100","0100","0101","0101","1000","1001","0111","0011","0011","0011","0101","1000","0110","0110","0110","0100","0011","0100","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","1000","0111"),
("0101","0100","0110","0110","0110","0110","0101","0101","0010","0010","0010","0011","0011","0010","0010","0010","0011","0010","0010","0011","0111","0100","0010","0010","0010","0001","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0010","0011","0011","0011","0011","0011","0010","0001","0001","0100","1010","1010","1011","0101","0010","0010","0001","0001","0010","0011","0101","0100","0100","0101","0101","0101","0101","0101","0011","0001","0010","0100","0101","0100","0100","0100","0100","0001","0010","0010","0111","1100","1100","1100","1100","1100","1100","1100","1100","1011","1100","1100","0100","0010","0011","0011","0010","0001","0010","0100","0100","0100","0100","1011","1101","1101","1101","1101","1101","1011","1000","0110","0111","0111","0111","0111","0111","0111","0110","0101","0100","0011","0010","0100","1001","1001","1000","1000","0110","0100","0011","0011","0011","0011","0100","0100","0011","0100","0011","0011","0011","0110","0110","0110","0110","0110","0110","0110","0100","0100","0101","0011","0010","0101","0100","0011","0011","0100","0011","0100","0100","0110","0101","0101","0010","0001","0001","0011","0010","0001","0001","0001","0001","0001","0001","0010","0001","0010","0100","0011","0010","0010","0001","0001","0001","0010","0010","0010","0100","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0110","1000","1001","1001","1010","1010","1011","1011","1011","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1011","1010","1010","1001","0111","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0101","0101","0010","0010","0010","0010","0010","0010","0110","1000","0110","0101","0101","0101","0101","0110","0111","0111","0111","0110","0101","0100","0001","0001","0001","0011","0111","0111","0111","0110","0110","0110","0110","0101","0110","0110","0110","0111","1000","0111","0111","0110","0100","0001","0010","0010","0011","0101","0101","0111","0110","0110","0110","0101","0100","0100","0101","0101","0110","0101","0100","0100","0100","0100","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0100","0111","1001","1000","1001","0101","0100","0111","0111","1000","1000","0110","0101","1000","0110","0110","1000","0110","0110","0100","0101","0101","0011","0010","0110","0110","0101","0010","0010","0010","0011","0111","1000","0111","0011","0010","0010","0010","0010","0010","0010","0011","1010","0111","0111","0111","0010","0001","0101","0100","0111","0100","0001","0101","0101","0100","0110","0110","0110","0101","0011","0010","0011","0011","0100","0110","0101","0110","0110","0101","0100","0010","0011","0011","0010","0100","0101","0110","0101","0101","0110","0100","0010","0010","0010","0011","0100","0101","0101","0101","0100","1000","1001","1010","0101","0011","0011","1000","1010","1001","1001","1001","1010","1000","1001","0111","1000","1001","1010","1001","1000","0110","0111","0100","0010","0010","0110","0111","0110","0101","0110","0111","0100","0100","0101","0111","0110","0110","0100","0110","0101","0100","0100","0101","1000","1000","0111","0100","0011","0011","0011","0011","0011","0011","0011","0011","0101","1001","0111","0010","0010","0001","0011","1000","0111","0101","0100","0011","0100","0011","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0001","0100","0110"),
("0100","0010","0010","0011","0101","0110","0101","0100","0010","0010","0010","0011","0100","0101","0101","0110","0110","0100","0011","0101","1000","0111","0011","0010","0010","0011","1000","1000","1000","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0010","0011","0011","0011","0100","0101","0101","0101","0101","0011","0011","0011","0100","0101","0110","0101","0101","0011","0011","0011","0011","0011","0100","0100","0101","0101","0100","0100","0100","0011","0011","0011","0011","0001","0001","0001","0000","0101","1001","1000","1000","0111","0100","0101","0110","1011","1011","1011","1001","0111","1000","1000","1010","1000","0110","0101","0011","0011","0011","0011","0100","0110","0110","0110","0110","1010","1100","1011","1100","1101","1100","1101","1101","1101","1101","1100","1011","1011","1100","1100","1011","0100","0011","0011","0011","0011","0100","0101","0110","0110","0101","0011","0100","0111","0101","0110","0111","0111","0110","0111","0110","0110","0111","0111","0111","0111","1000","0111","1000","0110","0010","0011","0100","0010","0001","0011","0011","0010","0010","0010","0010","0010","0011","0100","0101","0101","0011","0001","0010","0100","0011","0001","0001","0001","0001","0001","0010","0001","0001","0010","0101","0101","0100","0011","0010","0001","0010","0011","0011","0101","0011","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0101","1011","1011","1011","1011","1011","1100","1100","1100","1100","1011","1100","1100","1100","1100","1100","1100","1100","1100","1100","1011","1010","1010","1011","1011","1000","0100","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0010","0010","0001","0010","0010","0110","1000","0110","0101","0101","0101","0101","0110","0111","0111","1000","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0110","0101","0101","0101","0110","0110","0111","0111","1000","1000","0111","0110","0110","0110","0111","0111","0111","0111","0110","0110","0110","0110","0110","0101","0100","0100","0101","0101","0110","0110","0100","0100","0100","0101","0011","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0110","1001","0111","1000","0111","0101","0100","1000","0110","1000","0101","1001","1000","1000","0111","1000","1000","0111","0111","0110","0010","0100","0110","0110","0011","0010","0010","0011","0110","0111","0110","0100","0011","0010","0010","0010","0010","0010","0010","0100","0111","1000","0011","1000","0001","0001","0101","0100","0111","0100","0001","0100","0101","0100","1000","1000","0110","0101","0011","0010","0011","0011","0100","0110","0111","1000","1000","0111","0101","0011","0011","0011","0011","0101","0111","1000","0111","0110","0110","0101","0010","0011","0011","0011","0101","0110","0111","0111","0101","1000","1001","1010","0110","0011","0011","1000","1010","1001","1001","1001","1010","1000","1000","0011","0111","0111","1010","1001","1000","0110","0111","0100","0011","0011","0110","0111","0110","0101","0110","0111","0011","0100","0011","0111","0111","0110","0101","0111","0101","0011","0100","0100","1000","1000","0111","0010","0001","0001","0001","0001","0001","0001","0001","0001","0101","1001","0111","0101","0101","0001","0010","0101","0101","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0010","0001","0100"),
("0101","0010","0001","0001","0010","0010","0010","0100","0110","0110","0110","0111","0111","0111","0111","0111","0111","0100","0110","1000","1010","1010","0101","0010","0010","0100","1000","1001","1000","0011","0010","0011","0100","0100","0011","0011","0011","0010","0011","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0011","0010","0010","0010","0100","0101","0110","0110","0110","0101","0011","0011","0010","0011","0101","0101","0110","0110","0011","0011","0011","0010","0011","0101","0110","0110","0110","0110","0110","0110","0101","0100","0011","0011","0010","0010","0010","0010","0101","1010","1010","1010","1000","0011","0010","0100","1011","1011","1100","1000","0001","0001","0010","1001","0100","0010","0011","0100","0100","0101","1000","0110","1001","0011","0010","0111","0111","1001","1011","1100","1110","1100","1011","1100","1100","1100","0101","0010","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0101","0110","0100","0100","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0011","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0011","0010","0010","0011","0011","0010","0010","0010","0100","0010","0001","0010","0111","1000","1000","0110","0010","0001","0010","0101","0111","1000","0101","0001","0010","0011","0010","0011","0010","0101","0100","0011","0110","0110","1010","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1100","1100","1100","1100","1100","1100","1011","1011","1011","1011","1010","1010","1010","1001","0101","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0011","0011","0011","0010","0110","1000","0110","0100","0101","0100","0101","0110","0110","0111","0111","0111","0110","0110","0110","0110","0111","0111","1000","1000","1000","0111","0111","0110","0101","0101","0110","0110","0111","1000","1000","1000","0111","0111","0101","0101","0101","0101","0101","0101","0101","0110","0111","0110","0110","0101","0101","0100","0101","0101","0110","0110","0100","0100","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0010","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0100","1000","1000","1001","0101","0101","0101","0111","0111","1001","0111","0111","0111","0110","0111","0110","0101","0111","0111","0101","0111","0101","0100","0010","0010","0011","0110","0110","0101","0100","0010","0100","0010","0010","0010","0010","0010","0011","0101","1000","1010","0110","1010","0110","0100","0101","0101","0101","0011","0010","0011","0100","0100","1000","0111","0110","0101","0011","0010","0011","0100","0100","0110","0110","1000","1001","0110","0101","0011","0011","0010","0100","0100","0111","1001","1000","0111","0110","0101","0010","0011","0011","0011","0101","0110","0111","1001","0101","1000","1001","1010","0110","0100","0011","1000","1001","1001","1001","1001","1001","1000","0111","0011","0110","0110","1001","1001","1000","0110","0111","0101","0011","0100","0110","0111","0110","0101","0110","0111","0011","0100","0011","0111","0111","0110","0101","0111","0110","0010","0011","0100","1000","1000","0111","0011","0010","0010","0010","0010","0010","0010","0010","0010","0101","1000","0110","0100","0110","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0011","0011","0011","0011","0001"),
("0111","0010","0001","0001","0001","0010","0010","0110","1000","1000","1000","1000","1000","1000","1000","1000","1000","0100","0110","1000","1001","1000","0111","0100","0100","0100","0111","1001","0111","0010","0010","0011","0100","0100","0011","0011","0011","0011","0100","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0011","0011","0011","0010","0100","0101","0110","0101","0101","0101","0100","0011","0010","0100","0101","0101","0110","0101","0011","0011","0100","0011","0100","0101","0110","0110","0110","0110","0110","0110","0101","0100","0011","0011","0010","0100","0100","0101","0100","1000","1010","1010","1001","0011","0010","0011","0101","0110","0111","0101","0011","0010","0010","0101","0011","0010","0010","0100","0101","0110","0111","0110","0111","0011","0010","0101","0110","0111","1000","1001","1001","1001","1000","1001","1000","1001","0100","0010","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0010","0001","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0011","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0100","1010","0110","0011","0011","1000","0110","0011","0101","0101","0111","0100","0010","0100","1010","1010","1001","1001","0100","0010","0011","1001","1001","1010","1000","0011","0101","0101","0100","0100","0011","0111","0110","0100","0110","0111","1001","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1100","1100","1011","1010","1011","1011","1011","1100","1011","1011","1010","1010","1011","1010","0110","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","1001","1000","0100","0011","0100","0100","0100","0100","0100","0110","1000","0101","0100","0101","0101","0101","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0111","1000","1000","1000","0111","0111","0110","0101","0101","0101","0110","0111","1000","1000","1000","0111","0111","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0110","0101","0101","0100","0101","0101","0110","0110","0100","0100","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0110","1000","1000","1000","0111","0100","1000","1001","1001","0111","0111","0111","1001","0110","0110","0101","0101","0101","0111","1000","0110","0010","0001","0100","0111","0111","0100","0010","0100","0011","0100","0011","0010","0010","0010","0010","0011","0110","0111","1000","0111","0111","0110","0011","0011","0011","0011","0011","0010","0011","0011","0100","1000","0111","0110","0101","0100","0011","0100","0101","0100","0110","0110","0111","1000","0101","0100","0011","0011","0010","0011","0100","0110","1001","1000","0111","0110","0101","0011","0011","0100","0100","0101","0110","1000","1001","0101","1000","1001","1010","0110","0100","0100","1000","1001","1001","1001","1000","1001","0111","0111","0011","0110","0110","1000","1000","1000","0110","0111","0101","0011","0100","0110","0111","0111","0110","0110","0111","0011","0100","0100","0111","0111","0110","0101","0111","0101","0011","0100","0100","1000","1000","0101","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100"),
("0111","0011","0010","0010","0010","0011","0011","0110","1000","1000","1000","1000","1001","1001","1001","1001","1001","0100","0110","1000","1001","1001","1000","0111","0111","0111","0110","1000","0100","0010","0010","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0011","0011","0101","0101","0101","0110","0101","0100","0100","0100","0100","0101","0101","0110","0110","0110","0111","0111","0111","0111","0110","0101","0101","0110","0111","0101","0110","0100","0110","1001","1010","1001","0011","0010","0010","0011","0100","0101","0100","0011","0010","0010","0010","0010","0010","0010","0100","0101","0110","0110","0110","0101","0011","0010","0011","0101","0101","0101","0110","0110","0110","0110","0110","0110","0101","0011","0010","0010","0010","0001","0001","0011","0101","0101","0101","0101","0110","0100","0011","0011","0011","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0001","0010","0011","1000","0101","0010","0011","0110","0101","0010","0010","0101","0101","0110","1011","0110","0111","0101","1010","1000","0100","0110","0110","1000","0101","0011","1000","1011","1010","1010","1011","1000","0100","0110","1011","1001","1011","1010","0110","0111","0110","0100","0101","0100","0111","0101","0111","0111","1001","1000","1011","1011","1001","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1010","1010","1011","1011","0111","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0010","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0011","0011","0011","0100","0011","0100","0101","0100","1000","1000","0100","0010","0011","0011","0100","0100","0100","0111","1001","0110","0101","0101","0101","0101","0101","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","0110","0110","0101","0110","0110","0111","0111","1000","1000","1000","0111","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0101","0101","0101","0101","0101","0111","0110","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0011","0010","0011","0011","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0100","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0100","0110","0111","1000","1000","1000","0101","1000","0111","1000","1000","0101","1010","0011","1000","0101","0101","0100","0110","0111","0100","0100","0100","0111","0111","0011","0010","0010","0011","0101","0011","0101","0010","0010","0011","0100","0110","0111","0011","0101","0101","0010","0010","0011","0100","0011","0010","0010","0001","0100","0101","0100","0110","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0110","0101","0101","0010","0100","0101","0101","0100","0101","1000","0111","0111","0111","0101","0101","0101","0101","0101","0101","0110","0111","1000","0101","0111","1001","1000","0110","0110","0101","0111","1001","1001","0111","0100","0100","0100","0101","0100","0100","0100","0101","0101","0111","0110","0110","0100","0100","0100","0101","0111","0110","0101","0110","0101","0100","0100","0100","0110","0111","0110","0101","0110","0100","0100","0100","0100","0111","0110","0100","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100"),
("1000","0100","0010","0010","0011","0011","0011","0101","0111","0111","0111","1000","1000","1010","1010","1001","1001","0110","0111","1000","1001","1000","1001","0111","0101","0100","0100","0100","0011","0011","0010","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0110","0110","0101","0101","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0100","0101","0101","0101","0110","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0110","0101","0100","0100","0011","0011","0011","0010","0001","0001","0001","0011","0101","0011","0100","1001","1010","1001","0101","0100","0011","0011","0101","0101","0100","0011","0010","0010","0011","0010","0010","0011","0101","0110","0110","0110","0110","0101","0011","0010","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0011","0010","0010","0010","0010","0100","0101","0100","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0100","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0011","0111","1001","0011","0010","0110","1001","0100","0010","0101","1010","0111","1010","1011","0110","1010","0110","1011","1001","0100","0101","0111","1001","0100","0100","1001","1100","1010","1010","1100","1000","0100","0110","1100","1010","1010","1011","1000","0111","0111","0101","0101","0100","0111","0111","0111","0111","1001","1000","1010","1000","0111","1000","1010","1011","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1100","1011","1011","1010","1011","1011","1011","1000","0011","0011","0011","0011","0011","0100","0100","0100","0101","0110","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0100","0011","0100","0101","0100","0011","0011","0010","0010","0011","0011","0011","0011","1000","1001","0111","0101","0101","0101","0101","0110","0110","0111","0111","1000","1000","0111","0111","1000","1000","0111","0111","1000","1001","1000","0111","0111","0110","0110","0111","0110","1000","1000","1000","1000","1000","0111","0110","0111","0110","0110","0110","0111","0111","0110","0110","0110","0110","0101","0101","0101","0101","0101","0110","0110","0011","0100","0100","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0101","0011","0011","0010","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0011","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","0100","0011","0110","1000","1010","1000","0101","0111","0111","1001","0110","1000","0011","0111","0100","0110","0110","0101","0110","0101","0111","0111","0101","0011","0010","0010","0010","0010","0101","0011","0101","0100","0110","1000","0111","0101","0011","0001","0100","0111","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0111","0110","0110","0110","0110","0101","0101","0101","0110","0101","0110","0110","0110","0110","0111","0101","0111","0111","0110","0100","0100","0110","0110","0110","0110","0111","0110","0101","0101","0110","0110","0110","0111","1000","0101","1000","1010","1001","1010","1001","1001","1001","1001","1001","1000","0111","0110","0101","0110","0110","0110","0111","0111","0111","1000","0110","0111","1000","0111","0111","1000","0111","0111","0110","0110","1000","0111","0111","0111","0111","0111","0111","0101","0111","0111","0111","0111","0111","0111","0100","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011"),
("1001","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","1000","1000","1000","0110","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0100","0101","0101","0101","0101","0101","0101","0101","0110","0101","0011","0010","0011","0011","0011","0100","0100","0101","0110","0110","0110","0110","0101","0101","0110","0101","0110","0101","0100","0011","0011","0011","0010","0100","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0101","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0101","1001","1010","1001","1000","1001","1000","0011","0101","0110","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0011","0011","0011","0100","0101","0101","0100","0100","0100","0100","0100","0011","0011","0100","0100","0010","0010","0101","1001","1001","0110","0100","0110","0111","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0100","0100","0011","0010","0011","0011","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0011","0010","0010","0100","0100","0010","0011","0110","0101","0110","1011","1010","0111","1010","0111","1011","0111","0101","0101","1000","1000","0101","0101","1010","1100","1001","1001","1011","1000","0101","0101","1011","1010","1010","1010","1010","0111","0111","0110","0101","0100","0100","0100","0101","0111","0111","0111","0111","1001","0011","0111","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1001","0101","0011","0011","0011","0100","0100","0100","0100","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0100","0011","0100","0101","0100","0011","0011","0011","0011","0011","0011","0100","1000","1001","0111","0101","0101","0101","0101","0110","0110","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","1001","1001","1000","0111","0111","0111","0110","0110","0110","0111","1000","1000","1000","0111","0111","0110","0110","0110","0110","0110","0110","0111","0110","0111","0110","0110","0110","0101","0101","0101","0101","0111","0111","0100","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0010","0010","0010","0010","0011","0100","0100","0011","0100","0101","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","0101","0101","0100","0011","0110","1000","1000","0111","0111","0101","1001","1001","1000","0110","0111","0110","0111","0100","0100","0011","0111","1000","0110","0011","0010","0010","0010","0010","0010","0101","0111","1000","0111","0101","0100","0011","0010","0010","0010","0100","1000","0011","0011","0011","0010","0010","0100","0100","0100","0011","0011","0100","0111","0110","0100","0100","0100","0101","0110","0101","0011","0100","0101","0110","0101","0101","0101","0101","0101","0101","0101","0011","0100","0110","0110","0110","0101","0100","0101","0101","0101","0101","0100","0101","0111","1000","0101","1000","1010","1001","1010","1001","1010","1010","1001","1001","1000","0111","0110","0111","1000","1000","1000","1000","1000","1000","1000","0110","0111","0110","0101","0110","1000","1000","0111","0110","0110","1000","0110","0110","0111","1000","0111","0110","0101","0111","0111","0110","0110","0111","1000","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011"),
("1000","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0110","0110","0100","0001","0000","0000","0000","0000","0001","0011","0011","0011","0011","0011","0011","0011","0011","0010","0100","0101","0101","0101","0101","0101","0110","0101","0010","0010","0010","0010","0010","0101","0110","0100","0011","0101","0110","0110","0110","0101","0110","0101","0101","0101","0110","1001","1010","0111","1000","1000","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0101","0101","0100","0010","0010","0010","0010","0100","0100","0100","0110","0110","0110","1000","0110","0111","1000","1001","0110","0010","0010","0010","0011","0100","0011","0010","0011","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0101","1001","1001","1001","1001","0110","0100","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0100","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0011","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0111","1011","1010","1000","1010","1000","1011","0111","0010","0101","1000","0110","0100","0110","1011","1011","1001","1000","1011","1001","0101","0101","1010","1011","1001","1011","1010","0111","0110","0110","0101","0100","0100","0100","0101","0111","0110","1000","0101","1000","1000","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1001","0101","0011","0011","0011","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0100","0110","0100","0011","0100","0101","0101","0101","0101","1000","1010","1010","1000","0110","0101","0101","0110","0111","0111","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","1010","1010","1000","1000","1000","0111","0111","0111","0110","0111","1000","1001","1001","1001","1001","1000","0111","0111","0111","0110","0110","0110","0110","0110","0110","0101","0100","0100","0100","0100","0100","0101","0101","0100","0010","0000","0000","0001","0001","0001","0010","0010","0010","0001","0010","0001","0010","0110","0111","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0011","0010","0010","0011","0011","0011","0100","0010","0010","0010","0011","0011","0100","0110","0011","0011","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0110","0100","1000","0110","0101","0011","0101","1000","0111","1000","1000","1001","1010","1000","0111","1000","0110","0111","0110","0100","0110","0111","0101","0011","0100","0010","0010","0011","0101","0110","0111","0110","0100","0100","0010","0010","0010","0010","0010","0101","0100","1000","0110","0110","0011","0010","0011","0101","0101","0011","0011","0011","0100","0111","0110","0101","0101","0101","0111","0111","0110","0101","0110","0110","0110","0101","0011","0010","0010","0010","0010","0011","0100","0100","0101","0110","0110","0101","0101","0101","0111","0111","0101","0100","0101","0111","1000","0101","1000","1010","1001","1010","1001","1010","1001","1001","1001","1000","1000","0110","0110","0110","0111","0110","1001","1000","1000","1000","0110","0110","0101","0110","0110","0110","0111","0111","0110","0110","0110","0101","0110","0101","0110","0111","0110","0101","0111","0101","0101","0101","0101","0110","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0001","0001","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0010"),
("0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0001","0001","0001","0001","0000","0001","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0011","0100","0100","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0110","1011","1100","1010","1010","1010","0111","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0100","0010","0011","0011","0101","0101","0100","0100","0011","0100","0100","0100","0101","0111","0110","0101","0110","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0111","1001","1001","1001","1001","1001","0110","0100","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0101","0100","0101","0100","0010","0010","0010","0010","0011","0110","0100","1000","1011","1001","1001","1000","1001","1100","1100","0110","0101","0111","0111","0111","1001","1010","1010","1000","1000","1011","1010","0111","0111","1001","1010","1000","1001","1010","1001","0110","0110","0110","0100","0101","1001","1000","0110","0110","0111","0111","0111","1001","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0101","0100","0010","0100","0110","0110","0111","0111","0110","0101","0110","0101","0100","0011","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0110","0110","0111","1000","1001","1000","1000","0111","0110","0101","0110","0110","0101","0101","0110","0111","0111","0111","0111","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0010","0010","0010","0011","0010","0010","0000","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0111","0111","0100","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0010","0001","0011","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0100","0010","0001","0010","0010","0010","0001","0010","0001","0010","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0001","0001","0010","0100","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0011","0100","0111","1001","1010","1000","0100","0011","0110","0111","1010","1010","1010","1001","1001","1000","0111","0110","0111","0111","0101","0011","0100","0011","0101","0101","0111","0111","0110","0011","0010","0100","0010","0100","0010","0001","0001","0001","0010","0011","0100","1001","0101","0101","0100","0010","0011","0011","0011","0011","0011","0011","0100","0111","0110","0110","0101","0100","0011","0011","0100","0101","0110","0110","0110","0101","0011","0010","0001","0010","0010","0010","0011","0100","0101","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0111","1000","0101","1000","1010","1001","1001","1000","1001","1001","1001","1001","1001","1000","0101","0101","0101","0101","0101","0101","1000","1000","1000","0110","0101","0110","0110","0110","0110","0110","0111","0110","0101","0110","0110","0110","0111","0110","0110","0110","0101","0110","0101","0110","0111","1010","0111","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0001","0001","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0010"),
("0100","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0001","0000","0001","0001","0000","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0100","0011","0011","0101","1011","1100","1011","1011","1011","0110","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0111","1001","1001","1001","1001","1001","0111","0100","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0100","0100","0011","0100","0100","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0100","0101","0100","0100","0100","0010","0010","0101","0111","0111","1001","0111","1001","1010","1000","1000","0111","1000","1001","1001","1001","0110","0110","1000","1000","0111","0111","0111","0111","1000","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1001","1001","1001","1001","1000","1000","1000","0111","1001","1000","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1001","0110","0100","0011","0011","0011","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0110","0100","0010","0011","0101","0110","0110","0110","0110","0101","0100","0011","0011","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0011","0011","0011","0100","0100","0010","0000","0000","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0111","0110","0100","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0100","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0001","0001","0001","0001","0001","0001","0000","0001","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0001","0010","0100","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0100","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0010","0010","0010","0011","0101","0100","0100","0100","0100","0110","1001","1001","0111","0101","0111","1000","1001","1001","1010","1001","1001","0111","0111","1000","0110","0010","0010","0101","0111","1000","0110","0011","0010","0001","0001","0010","0100","0010","0011","0001","0001","0001","0010","0010","0010","0010","1000","0101","0101","0110","0010","0010","0010","0010","0100","0011","0011","0100","0111","0110","0110","0101","0011","0010","0010","0011","0011","0110","0110","0110","0101","0101","0100","0010","0010","0010","0001","0100","0101","0110","0110","0110","0110","0101","0010","0010","0010","0010","0100","0110","0111","1000","0101","1000","1001","1001","0100","0011","0011","1000","1001","1000","1000","1000","0101","0010","0010","0011","0011","0101","1000","1000","1000","0110","0110","0011","0010","0010","0100","0111","0111","0110","0101","0101","0011","0011","0011","0101","0110","0110","0101","0101","1000","1010","1100","1011","0101","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0010","0001","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0011","0011","0011"),
("0100","0101","0101","0100","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0000","0000","0001","0001","0000","0001","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0110","0110","0110","0110","0110","0111","0110","0110","0101","0101","0100","0100","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0111","0111","0110","0110","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0110","1001","1001","1001","1001","1001","0111","0100","0101","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0011","0011","0101","0101","0101","0101","0101","0100","0010","0010","0101","0110","0101","0100","0100","0101","0010","0011","0010","0011","1000","1001","1001","1001","1000","1000","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","1000","1000","1000","1000","1000","0111","1000","1000","1001","1010","1010","1001","1001","1010","1010","1001","1001","1010","1001","1010","1001","1000","0111","1000","0111","0111","0111","0110","0100","0100","0101","1000","1010","1010","1010","1010","1011","1011","1011","1011","1011","1010","1010","1010","1001","1001","1001","1001","1000","1000","1000","0111","0111","0111","0111","0110","0110","0110","0101","0101","0101","0100","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0101","0110","0011","0011","0101","0101","0101","0110","1000","0111","0101","0100","0100","0011","0011","0100","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0101","0110","0111","0101","0101","0100","0011","0100","0101","0011","0011","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0011","0100","0100","0100","0101","0101","0011","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0110","0110","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0110","0010","0010","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0110","0011","0011","0011","0011","0010","0010","0001","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0011","0010","0001","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0011","0011","0111","0110","0011","0100","0100","0011","0100","0101","0110","1000","1001","1010","1000","1010","1001","1010","1001","0111","0110","0101","0100","0110","0110","0110","0101","0100","0011","0001","0001","0001","0010","0001","0100","0010","0011","0010","0001","0001","0001","0001","0001","0001","0111","0101","0100","0110","0010","0010","0011","0011","0011","0010","0011","0100","0110","0110","0110","0101","0011","0010","0010","0011","0100","0110","0110","0110","0110","0101","0101","0010","0010","0011","0010","0101","0110","0110","0110","0110","0110","0101","0011","0010","0011","0011","0101","0110","0111","1000","0101","1000","1010","1010","0100","0010","0010","1000","1001","1001","1000","1000","0101","0010","0010","0010","0010","0101","1000","1000","1000","0110","0110","0011","0011","0011","0100","0111","0111","0110","0110","0101","0010","0010","0001","0101","0110","0110","1000","1010","1011","1011","1001","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0101"),
("0100","0100","0101","0100","0101","0100","0110","0101","0011","0010","0010","0010","0011","0011","0011","0011","0011","0100","0100","0100","0101","0100","0100","0101","0100","0011","0011","0011","0011","0011","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0101","1000","1001","1001","1001","1001","0111","0100","0101","0110","0110","0110","0110","0110","0111","0111","0100","0011","0101","0101","0100","0100","0101","0110","0110","0101","0100","0011","0010","0010","0011","0011","0011","0100","0101","0100","0100","0100","0101","0100","0110","0111","0110","0101","0100","0100","0010","0010","0010","0010","0010","0100","0111","0110","0110","1000","1001","1001","1001","0101","0010","0011","0100","1001","1010","1010","1010","1010","1010","1000","1000","1001","1001","1001","0100","0011","0011","0111","0111","0100","0101","0100","0010","0010","0011","0011","0011","0100","0011","0100","0101","1000","0111","0111","0111","0111","0110","0110","0101","0101","0101","0101","0101","0101","0100","0011","0100","0011","0011","0011","0100","0101","0101","0101","0101","0101","0100","0010","0010","0001","0001","0001","0010","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0110","0110","0111","0011","0001","0011","0100","0100","0100","0111","1000","0110","0101","0100","0011","0100","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","1000","1001","0110","0110","0101","0011","0100","0101","0100","0100","0101","0110","0110","0110","0110","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0011","0100","0100","0100","0101","0110","0011","0000","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0110","0110","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","0101","0010","0001","0001","0001","0001","0010","0001","0001","0010","0001","0001","0001","0010","0001","0001","0001","0010","0101","0011","0100","0011","0011","0011","0010","0010","0011","0011","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","0100","0010","0100","0010","0010","0010","0011","0011","0011","0011","0100","0100","0101","0101","0110","0110","0101","0100","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0010","0101","0111","0011","0100","0100","0011","0100","0010","0010","0011","0110","1000","1000","1001","1010","1001","1000","0111","0110","0110","0101","0100","0010","0010","0100","0011","0100","0010","0010","0001","0001","0001","0011","0011","0011","0010","0001","0001","0001","0001","0001","0001","0110","0101","0100","0111","0001","0010","0011","0011","0010","0011","0100","0100","0110","0110","0110","0101","0011","0010","0010","0011","0011","0110","0110","0101","0101","0101","0110","0010","0011","0010","0011","0101","0110","0110","0101","0110","0110","0101","0010","0010","0011","0011","0100","0110","0111","1000","0101","1000","1010","1010","0101","0010","0010","1000","1001","1001","1001","1000","0101","0010","0010","0010","0010","0101","1001","1000","1000","0110","0110","0100","0101","0101","0101","0111","0111","0110","0101","0101","0101","0110","0101","0110","1000","1010","1011","1011","1011","1001","0110","0111","0111","0110","0111","0111","0110","0000","0010","0111","0111","0111","0110","0111","0111","0100","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0100","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0101"),
("0100","0100","0101","0101","0100","0011","0100","0011","0010","0001","0001","0010","0010","0010","0011","0011","0011","0100","0110","0110","0111","0111","0110","0110","0100","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0010","0100","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0011","0011","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0101","1000","1001","1001","1001","1001","1000","0100","0101","0110","0110","0110","0101","0100","0100","0001","0011","0101","0101","0100","0100","0101","0110","0110","0101","0100","0100","0010","0010","0011","0011","0110","1000","1000","1000","1001","1001","1010","1010","1001","1001","0110","0011","0010","0010","0011","0011","0011","0011","0011","0111","1001","0111","0111","1000","1010","1010","1010","0110","0011","0011","0100","1001","1010","1011","1011","1011","1010","1001","1001","1010","1010","1010","0011","0010","0011","1001","0111","0011","0100","0011","0100","0011","0010","0011","0011","0010","0011","0010","0100","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0011","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0101","0111","0011","0010","0011","0011","0011","0011","0111","1000","0110","0101","0100","0100","0100","0101","0110","0110","0111","0111","0110","0111","0110","0111","0110","0110","0111","1000","1000","0110","0110","0101","0100","0100","0101","0100","0101","0110","0111","0110","0110","0110","0100","0101","0101","0101","0110","0101","0110","0110","0110","0110","0101","0101","0100","0100","0100","0100","0101","0101","0011","0000","0001","0001","0010","0010","0011","0011","0011","0010","0011","0100","0011","0100","0110","0110","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0011","0011","0010","0010","0011","0010","0011","0100","0100","0011","0011","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0110","0100","0101","0001","0001","0001","0001","0010","0101","0101","0100","0011","0011","0011","0100","0011","0100","0100","0100","0100","0100","0101","0100","0011","0110","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0110","0110","0111","0110","0101","0011","0101","0100","0101","0110","0111","0111","0110","0110","0111","0111","0111","0111","1000","0110","0101","0101","0011","0011","0100","0100","0100","1000","0111","0111","0111","0111","0110","0110","0110","0111","1001","1010","1001","0111","0111","0110","0101","0101","0101","0101","0101","0110","0101","0101","0100","0100","0011","0010","0010","0011","0011","0011","0011","0001","0001","0001","0001","0001","0001","0101","0110","0100","0111","0010","0010","0010","0010","0010","0011","0011","0011","0101","0101","0110","0101","0011","0010","0010","0100","0011","0110","0110","0100","0011","0100","0110","0011","0011","0001","0011","0100","0100","0011","0101","0110","0110","0101","0010","0010","0011","0011","0100","0110","0111","1000","0101","1000","1001","1010","0101","0010","0010","1000","1001","1001","1000","1000","0110","0010","0011","0001","0011","0101","0111","1000","1000","0110","0110","0100","0101","0011","0100","0111","0111","0110","0110","0101","0011","0110","1000","1010","1011","1011","1011","1011","1011","1010","0111","1000","1000","1000","1000","1000","0111","0100","0101","1000","1000","1000","0111","1000","1000","0101","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0101","0111","0111","0111"),
("0101","0101","0101","0100","0101","0101","0100","0010","0011","0010","0010","0010","0100","0100","0011","0011","0100","0110","0101","0101","0101","0100","0101","0110","0110","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0011","0011","0011","0100","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0100","0011","0011","0011","0100","0100","0011","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0101","1000","1001","1001","1001","1001","1000","0100","0101","0110","0110","0110","0100","0011","0010","0100","0101","0101","0101","0101","0100","1000","1010","1001","1001","1001","0011","0011","0011","0010","0110","0111","0111","1000","1001","1001","1001","1000","1001","0111","0101","0011","0011","0101","0011","0010","0010","0010","0010","0101","1000","1001","1001","1001","1001","1010","1001","0110","0010","0010","0100","1000","1001","1001","1001","1001","1001","1001","1000","1001","1001","1000","0011","0010","0011","0111","0110","0101","0101","0100","0101","0100","0100","0011","0010","0010","0010","0010","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0101","0101","0101","0101","0101","0100","0010","0010","0100","0101","0101","0101","0101","0110","0110","0110","0101","0111","0110","0110","0101","0101","0101","0100","0100","0100","0100","0011","0011","0111","0101","0011","0100","0010","0011","0011","0011","0010","0011","0110","0111","0110","0100","0100","0100","0101","0110","0111","0111","1000","1000","1000","1000","1000","1001","1000","1000","1000","0111","0111","0110","0101","0101","0100","0100","0101","0100","0101","0110","0110","0111","0110","0101","0110","0110","0101","0110","0111","0110","0110","0111","0110","0110","0101","0101","0100","0100","0100","0101","0101","0110","0011","0000","0001","0010","0011","0100","0100","0100","0100","0100","0101","0101","0101","0101","0110","0110","0100","0100","0110","0110","0110","0110","0110","0110","0110","0101","0110","0101","0110","0101","0101","0110","0101","0101","0110","0101","0100","0010","0100","0111","0111","0110","0111","0111","1000","0110","0101","0110","0111","0110","0111","0110","0110","0110","0111","0101","0101","0011","0011","0011","0011","0010","0101","0101","0101","0101","0110","0110","0110","0101","0101","0101","0101","0101","0101","0110","0100","0011","0101","0110","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0011","0011","0101","0100","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0100","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0101","0110","1010","1001","0111","0111","0111","0111","0110","0101","0101","0101","0101","0110","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0101","0110","1001","1001","1001","1010","0101","0001","0010","0011","0011","0100","0011","0011","0110","0101","0101","0101","0100","0011","0011","0100","0100","0110","0101","0011","0010","0100","0101","0011","0100","0011","0100","0011","0011","0010","0101","0110","0110","0101","0011","0011","0011","0100","0100","0110","0111","0111","0101","0111","1001","1010","0101","0011","0011","1000","1001","0111","0111","0111","0110","0010","0011","0001","0011","0100","0110","0111","0111","0110","0101","0101","0101","0100","0100","0110","0110","0101","0101","0110","1001","1011","1011","1011","1011","1011","1011","1011","1011","1010","0111","1000","0111","0111","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","0111","0100","0010","0010","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0101","1000","0111","0111"),
("0101","0110","0101","0011","0100","0101","0011","0010","0100","0100","0101","0101","0101","0110","0011","0100","1000","1010","1010","1010","1001","1010","1001","1001","1010","1000","0100","0011","0011","0011","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0100","1000","1001","1001","1001","1001","1000","0101","0101","0110","0110","0110","0101","0011","0100","0101","0110","0101","0101","0101","0101","1000","1010","1010","1001","0011","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0010","0010","0010","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0011","0011","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0010","0011","0011","0100","0110","0101","0100","0100","0100","0100","0010","0011","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0110","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","1000","0110","0101","0101","0100","0100","0101","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0110","0101","0101","0100","0101","0101","0101","0101","0110","0111","0111","0111","0110","0101","0101","0101","0101","0110","0110","0110","0111","0111","0101","0101","0101","0100","0100","0100","0101","0110","0101","0011","0001","0001","0011","0011","0100","0100","0100","0101","0110","0110","0101","0101","0110","0111","0110","0100","0100","0101","0110","0110","0110","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0100","0010","0011","0111","0111","0111","1000","0111","0111","0111","0110","0111","0111","0111","1000","1000","0111","0111","0111","0101","0101","0100","0101","0101","0100","0100","0101","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0100","0100","0101","0101","0110","0110","0111","0111","0111","0111","0111","0110","0110","0110","0101","0100","0011","0011","0100","0100","0110","0111","0111","0111","1000","0110","0110","0111","0111","0110","0110","0101","0100","0011","0100","0100","0101","0100","0011","0011","0011","0010","0011","0101","0111","0110","1001","1011","1010","1001","0111","0111","1000","1001","1000","0101","0011","0001","0011","0010","0011","0010","0010","0010","0010","0001","0010","0011","0011","0011","0010","0011","0011","0011","0100","0100","0101","0110","0011","0100","0010","0001","0001","0010","0010","0011","0011","0011","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0101","0010","0100","0101","0110","0101","0110","0110","0101","0011","0010","0011","0101","0110","0110","0110","0101","0110","0110","0110","0110","0110","0111","1000","0101","0110","1000","1000","0101","0101","0101","0111","0111","0011","0011","0011","0101","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0101","0110","1001","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0111","0111","0111","0110","0110","0110","0101","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0100","0110","0110","0110"),
("0010","0011","0011","0100","0100","0011","0011","0011","0101","0111","0111","0110","0111","0101","0011","0110","1001","1010","1010","1001","1010","1011","1010","1001","1001","1001","0110","0011","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0101","1000","1001","1001","1001","1001","1001","0101","0101","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","0011","0100","1000","1011","1010","0101","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0010","0011","0011","0011","0100","0110","0111","0111","1000","0111","0110","0011","0100","0100","0100","0100","0101","0101","0101","0100","0100","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0100","0110","0110","0010","0011","0011","0100","0011","0011","0011","0011","0011","0011","0110","0111","0101","0101","0100","0100","0100","0110","0110","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0101","0101","0110","0101","0101","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0101","0101","0100","0100","0101","0101","0110","0110","0011","0001","0010","0010","0011","0100","0100","0101","0100","0110","0101","0101","0100","0101","0101","0101","0100","0100","0100","0101","0110","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0110","0110","0110","0101","0101","0011","0100","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0110","0110","0101","0101","0110","0101","0101","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0101","0101","0100","0100","0101","0110","0110","0101","0110","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0101","0100","0100","0101","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0101","0100","0011","0100","0100","0101","0100","0011","0101","0111","0111","0110","0101","0100","0111","1011","0111","0110","1010","1000","1000","1000","1001","1000","1000","0111","0111","0101","0011","0011","0010","0010","0010","0010","0010","0011","0010","0011","0010","0001","0001","0001","0001","0001","0001","0100","0101","0001","0010","0001","0001","0001","0001","0001","0001","0001","0011","0110","0101","0101","0110","0111","0111","0111","0111","0111","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0010","0010","0100","0101","0110","0110","0111","1000","1000","0111","1000","0111","0110","0111","0111","0101","0110","0110","0111","0111","0110","0110","0110","0101","0100","0100","0011","0011","0011","0100","0101","0011","0100","0011","0100","0011","0010","0011","0011","0011","0011","0101","0111","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1000","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0100","0100"),
("0010","0010","0011","0010","0010","0010","0011","0011","0011","0100","0011","0100","0100","0011","0011","1000","1001","1001","1000","1000","1010","1011","1001","1001","1000","1000","0110","0011","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0011","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0100","0011","0011","0100","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0111","1001","1001","1001","1001","1001","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","1000","0111","0011","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0010","0010","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0101","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0111","1000","1000","1000","0111","0111","0111","1000","1000","0111","0011","0100","0100","0100","0101","0101","0101","0101","0100","0101","0100","0110","0101","0100","0011","0101","0100","0010","0101","0101","0010","0110","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0111","0110","0101","0100","0100","0101","0110","0101","0110","0111","0111","0111","0111","0101","0111","0111","0111","0111","0111","0111","0110","0110","0110","0101","0101","0110","0101","0101","0110","0110","0111","0111","0111","0101","0110","0110","0101","0011","0101","0110","0110","0101","0101","0100","0100","0100","0100","0100","0101","0110","0101","0100","0001","0001","0010","0100","0100","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0100","0100","0101","0110","0110","0110","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0111","0110","0110","0101","0110","0100","0011","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0101","0101","0110","0110","0101","0101","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0100","0101","0110","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0110","0110","0110","0101","0011","0100","0101","0111","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0100","0011","0100","0100","0101","0101","0111","1000","0110","0101","0001","0100","0110","1010","1001","0100","0101","0111","1011","0111","1000","1001","0111","0101","0101","1000","1010","1000","0110","0011","0010","0010","0010","0010","0100","0010","0011","0001","0001","0001","0001","0001","0001","0001","0110","0101","0001","0010","0010","0001","0001","0001","0010","0010","0010","0011","0101","0101","0101","0101","0110","0111","0110","0111","0110","0110","0101","0101","0011","0011","0100","0100","0100","0011","0100","0010","0010","0100","0101","0101","0101","0111","1000","0111","0110","0110","0110","0101","0110","0111","0101","0111","1001","1000","1000","1000","1000","1000","0111","0110","0110","0101","0101","0101","0101","0110","0101","0110","0110","0110","0101","0101","0011","0011","0010","0100","1001","1011","1011","1010","1011","1011","1011","1010","1011","1011","1010","1010","1010","1010","1000","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011"),
("0010","0011","0011","0010","0010","0010","0010","0011","0101","0101","0101","0101","0010","0010","0100","1000","1001","1000","1000","1000","1001","1010","1000","1000","0111","0111","0111","0100","0010","0010","0010","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0100","0011","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0101","1000","1001","1001","1001","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0011","0010","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0101","0100","0101","0100","0100","0100","0100","0100","0100","0110","1000","1010","1001","1001","1001","1001","0111","0011","0111","1000","0111","0011","0100","0100","0010","0010","0001","0010","0010","0011","0101","0101","0110","0110","0100","0010","0110","0101","0001","0100","0110","0110","0100","0100","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0111","0111","0110","0100","0101","0100","0100","0101","0110","0111","0111","0111","0111","0100","0010","0100","0111","0110","0110","0111","0111","0111","0110","0110","0101","0101","0101","0101","0101","0110","0110","0111","0111","0110","0101","0101","0101","0010","0010","0011","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0110","0110","0101","0001","0010","0010","0011","0100","0100","0100","0100","0101","0101","0100","0100","0110","0101","0101","0100","0100","0101","0110","0110","0110","0111","0111","0111","0111","1000","0111","0111","0111","0110","1000","1000","0111","0111","0110","0110","0100","0011","0110","0111","1000","0111","0111","1000","0111","1000","0111","1000","1000","1000","1000","1000","0111","0111","0111","0101","0101","0110","0111","0101","0101","0110","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0110","0100","0100","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0101","0100","0100","0110","0111","0110","0110","0110","0111","0111","0111","0110","0110","0110","0110","0110","0101","0100","0011","0100","0100","0101","0101","0100","0101","0011","0100","0100","0101","0111","1010","0110","0101","0110","0101","1010","1010","0101","1001","1000","0110","0101","0011","0101","1000","1000","1000","0110","0100","0010","0001","0100","0010","0011","0001","0001","0001","0001","0001","0001","0011","1000","0101","0101","0101","0100","0010","0010","0001","0001","0010","0011","0011","0110","0110","0101","0101","0110","0110","0101","0111","0110","0101","0101","0100","0100","0010","0001","0010","0010","0010","0011","0100","0010","0100","0101","0101","0101","0110","0111","0111","0110","0110","0110","0101","0101","0110","0101","0110","0111","0111","0111","0111","0111","0110","0100","0011","0011","0011","0100","0100","0100","0100","0011","0011","0100","0011","0011","0011","0011","0100","0011","0011","0101","1010","1011","1011","0111","0100","0111","0110","0101","0111","1000","1001","1001","1001","1000","0101","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001"),
("0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0011","0011","0010","0010","0110","1001","1001","1000","1000","1001","1001","1010","1000","1000","0111","0111","1000","0101","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0011","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0111","1000","1001","1001","1001","1001","0111","0100","0100","0100","0100","0100","0101","0101","0100","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0011","0110","1000","1010","1001","1001","1001","1001","1001","1001","1000","0111","1000","0111","0100","0101","0101","0001","0001","0001","0001","0010","0010","0101","0110","0111","0110","0011","0001","0101","0100","0101","1000","0111","0100","0011","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0111","1000","0110","0101","0101","0100","0100","0101","0111","0111","0111","0111","0101","0011","0010","0001","0110","1000","0111","0111","0111","0111","0110","0110","0101","0101","0110","0101","0110","0110","0110","1000","0111","0110","0110","0110","0100","0001","0010","0011","0100","0101","0110","0110","0101","0101","0101","0100","0100","0100","0101","0101","0100","0010","0010","0011","0100","0100","0100","0100","0100","0101","0101","0100","0100","0110","0101","0101","0100","0100","0101","0110","0110","0110","0111","0110","0110","0111","0111","0110","0111","0111","0110","1000","1000","1000","1000","0110","0110","0100","0011","0110","0111","1000","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0101","0110","0111","0101","0101","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0110","0100","0100","0101","0110","0110","0110","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0101","0101","0100","0100","0101","0110","0110","0101","0110","0110","0101","0100","0110","0110","0110","0110","0110","0101","0100","0011","0100","0101","0101","0101","0010","0011","0100","0110","0111","0101","1010","0111","0110","0111","0110","0100","1000","1011","0111","0110","1010","0111","0111","0110","0011","0011","0011","0110","1001","1000","0110","0101","0100","0010","0011","0001","0001","0001","0001","0001","0001","0011","1000","0101","0101","0101","0011","0001","0001","0001","0001","0010","0010","0011","0101","0101","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0010","0001","0001","0010","0010","0010","0011","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0110","0111","1000","0111","0111","0111","0111","0101","0101","0100","0001","0010","0010","0010","0011","0011","0011","0100","0011","0010","0011","0101","0100","0101","0111","1010","1010","1010","0111","0011","1000","0111","0110","0110","0100","0101","0110","0110","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010"),
("0011","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0010","0010","0010","1000","1010","1010","0110","0111","1000","1001","1010","1000","1000","0110","0110","1001","0111","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0100","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0011","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0100","1000","1000","1001","1001","1001","1000","0101","0101","0101","0101","0101","0101","0101","0100","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0101","0101","0101","0101","0101","0101","0101","0101","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","1000","1001","1010","1001","1001","1001","1001","1001","1001","1001","1000","0111","0111","0101","0110","0101","0010","0010","0010","0010","0001","0010","0100","0101","0110","0101","0010","0001","0100","0011","0010","0111","0110","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0111","1000","0110","0101","0101","0100","0101","0110","0111","0111","0111","0111","0100","0011","0001","0001","0011","0111","0111","0111","1000","0110","0110","0110","0110","0101","0110","0101","0110","0110","0110","0111","0110","0110","0110","0110","0010","0001","0001","0011","0100","0110","0110","0101","0101","0101","0101","0100","0100","0101","0101","0101","0100","0001","0010","0010","0100","0100","0100","0101","0101","0101","0101","0101","0101","0110","0101","0101","0100","0100","0101","0110","0110","0111","0111","0110","0110","0111","0111","0110","0111","0110","0111","1001","1000","1001","1000","0101","0101","0011","0011","0110","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0110","0110","0101","0101","0111","0111","0101","0101","0110","0110","0110","0111","1000","1000","0111","0111","0111","0111","0111","1000","0111","0111","0101","0100","0100","0101","0101","0110","0111","0110","0111","0100","0100","0110","0111","0111","0110","0110","0110","0101","0101","0100","0100","0101","0110","0110","0101","0110","0101","0001","0001","0010","0110","0110","0110","0110","0101","0100","0011","0100","0100","0101","0101","0010","0011","0111","0111","0110","0110","1001","0101","0111","0110","0101","0100","0101","1001","1010","0011","1000","1010","1000","1000","0111","0010","0001","0010","0010","0101","0111","1001","1001","0110","0100","0001","0001","0001","0001","0001","0001","0010","1000","0100","0101","0011","0001","0001","0001","0001","0001","0010","0010","0010","0110","0101","0100","0100","0010","0001","0010","0010","0010","0100","0101","0101","0110","0100","0010","0001","0001","0010","0010","0010","0100","0110","0101","0101","0101","0100","0010","0010","0010","0010","0011","0100","0011","0100","0100","0100","0100","0110","0101","0100","0011","0011","0100","0100","0011","0100","0001","0001","0010","0010","0011","0011","0011","0101","0101","0100","0110","0110","0101","1000","1001","0111","0111","0110","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100"),
("0010","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0001","0001","0100","1001","1000","1000","0110","0110","1000","1001","1010","1001","1000","0110","0101","0111","0101","0011","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0100","0011","0011","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0100","0111","1000","1000","1000","0110","0101","0100","0101","0101","0101","0100","0100","0011","0011","0011","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0110","0101","0011","0100","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0011","0110","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0111","0101","0110","0100","0010","0010","0010","0010","0001","0010","0101","0101","0110","0101","0010","0010","0100","0011","0011","0110","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","1000","1000","0110","0101","0101","0101","0101","0110","0111","0111","0111","0110","0100","0010","0001","0001","0010","0110","0111","1000","1000","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0111","0110","0100","0001","0001","0001","0010","0100","0101","0110","0110","0101","0101","0100","0101","0101","0101","0101","0100","0100","0001","0001","0010","0011","0100","0100","0011","0100","0100","0101","0101","0101","0110","0101","0100","0100","0100","0101","0110","0111","0110","0110","0111","0111","0111","0110","0010","0100","0111","0110","1000","1001","1000","1000","0110","0101","0011","0011","0110","0111","0111","1000","0111","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0101","0101","0111","0110","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","1000","1000","0111","0110","0100","0100","0101","0101","0110","0110","0111","0100","0001","0001","0011","0111","0111","0110","0110","0110","0110","0101","0100","0100","0101","0110","0110","0110","0110","0011","0001","0001","0001","0100","0110","0110","0110","0110","0100","0011","0100","0100","0101","0100","0100","0110","0110","0110","0100","1010","0111","0110","0111","0100","0110","0011","0110","0101","1011","0111","0101","1010","1000","1000","0110","0111","0010","0001","0010","0001","0010","0100","0111","1001","0111","0110","0100","0001","0001","0001","0001","0010","1000","0010","0110","0010","0001","0001","0001","0001","0010","0001","0010","0010","0100","0101","0100","0100","0011","0010","0010","0010","0011","0101","0101","0101","0110","0100","0011","0010","0001","0010","0010","0011","0100","0110","0110","0111","0110","0101","0011","0010","0011","0010","0011","0101","0101","0100","0011","0011","0011","0101","0011","0010","0010","0000","0100","0011","0010","0100","0100","0101","0110","0111","0011","0010","0011","0101","0101","0100","0101","0101","0100","0100","0011","0011","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0100","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101"),
("0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0010","0110","0110","0100","0101","0100","0100","0111","1001","1001","1001","0111","0100","0100","0100","0100","0011","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0011","0011","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0111","1000","1000","1000","0110","0111","0110","0110","0110","0111","0101","0001","0001","0001","0001","0010","0010","0011","0100","0100","0100","0100","0100","0100","0110","0110","0011","0010","0010","0011","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0011","0111","1001","1001","1001","0111","1000","0111","0111","0111","0111","1000","1000","1000","1000","1000","0111","0101","0100","0001","0001","0010","0010","0001","0010","0100","0100","0101","0101","0010","0010","0100","0100","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","1000","1000","0110","0101","0101","0101","0101","0110","0111","0111","0111","0110","0100","0010","0001","0010","0001","0101","0111","0111","1000","0110","0110","0110","0110","0110","0110","0101","0110","0110","0111","0111","0111","0110","0110","0011","0001","0001","0001","0010","0100","0101","0110","0110","0110","0101","0100","0100","0101","0101","0101","0101","0101","0001","0001","0010","0011","0100","0011","0001","0010","0100","0100","0101","0101","0110","0101","0100","0100","0100","0101","0101","0110","0110","0110","0111","0110","0110","0011","0001","0001","0101","0110","0111","0110","0110","1000","0110","0110","0011","0011","0101","0111","0111","0111","0111","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0111","0110","0101","0101","0110","0110","0110","0101","0110","0110","0110","0110","0101","0111","0111","0111","0111","0110","0101","0100","0101","0101","0101","0110","0111","0101","0001","0001","0001","0001","0100","0111","0110","0110","0110","0110","0101","0100","0100","0101","0110","0110","0110","0101","0001","0000","0001","0001","0011","0110","0110","0110","0110","0100","0011","0100","0100","0110","0110","0111","0110","0011","0100","1000","1001","0111","1000","0110","0100","0110","0011","0110","0100","1000","1011","0110","1001","1001","0101","0111","0111","0111","0011","0001","0001","0001","0011","0010","0100","0110","1000","1001","0111","0101","0010","0001","0011","0111","0010","0111","0010","0001","0001","0001","0001","0001","0001","0001","0010","0100","0100","0100","0100","0011","0001","0010","0011","0010","0100","0101","0101","0101","0100","0011","0011","0100","0110","0111","1000","1001","0111","0110","0111","1000","1000","0110","0100","0011","0011","0011","0100","0100","0100","0011","0011","0010","0100","0100","0010","0010","0010","0111","1000","1000","1000","0111","0110","0110","0101","0100","0011","0100","0100","0011","0100","0011","0011","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101"),
("0011","0011","0011","0010","0011","0010","0010","0010","0001","0001","0001","0001","0011","1000","0111","0011","0011","0011","0011","0110","1000","0111","0111","0110","0011","0100","0011","0010","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0010","0110","0101","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0011","0110","1000","1000","0111","0101","0110","0101","0110","1000","1001","0111","0001","0001","0001","0001","0010","0010","0011","0100","0100","0100","0100","0100","0101","0101","0101","0100","0010","0010","0011","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0100","0100","0100","0100","0011","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0010","0101","1001","1001","1001","1000","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","1000","1000","0110","0101","0101","0101","0100","0101","0111","0111","0111","0110","0100","0010","0001","0010","0010","0100","1000","1000","1000","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110","0010","0001","0010","0001","0010","0100","0101","0110","0110","0110","0101","0100","0101","0101","0101","0101","0101","0101","0010","0010","0010","0011","0011","0001","0010","0001","0011","0101","0101","0101","0101","0101","0100","0100","0101","0110","0110","0110","0110","0110","0110","0111","0100","0001","0010","0001","0010","0101","0110","0101","0110","1000","0110","0101","0011","0011","0101","0110","0111","0111","0111","0110","0110","0110","0111","0111","0110","0110","0110","0101","0110","0111","0110","0101","0100","0101","0101","0100","0101","0110","0110","0110","0101","0101","0110","0110","0011","0001","0011","0101","0110","0110","0101","0101","0100","0100","0101","0101","0110","0111","0011","0001","0001","0001","0001","0010","0110","0110","0110","0110","0110","0101","0100","0101","0110","0110","0110","0110","0100","0001","0001","0001","0010","0010","0110","0110","0110","0110","0100","0011","0100","0101","0110","0110","0111","0010","0001","0101","1010","0111","0111","1000","0101","0100","0101","0011","0101","0101","0101","1010","1010","0111","1010","0111","0011","0111","0111","0111","0100","0001","0010","0011","0011","0011","0001","0010","0101","0111","0110","0101","0100","0101","0101","0011","0111","0001","0001","0001","0001","0010","0010","0001","0001","0010","0101","0101","0100","0100","0011","0001","0010","0011","0010","0100","0110","0101","0100","0100","0011","0011","0101","1000","1001","1010","1011","1011","1001","0110","0100","0101","0110","0100","0100","0100","0100","0100","0100","0101","0011","0001","0001","0100","0101","0011","0011","0100","0101","0101","0100","0011","0010","0010","0010","0010","0100","0100","0101","0101","0011","0100","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0101","0110","0110","0110","0101","0110","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0100","0101","0101","0101","0110","0110","0110","0110","0110","0110","0101","0101","0110","0110","0101","0101","0101","0110","0110","0110","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101"),
("0010","0010","0011","0010","0010","0010","0001","0001","0001","0001","0001","0001","0101","1001","1001","0010","0011","0100","0101","0101","0100","0100","0011","0100","0100","0101","0100","0001","0110","0110","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0010","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0100","0110","0110","0110","0100","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0110","0011","0010","0010","0010","0010","0010","0100","0111","1000","0111","0011","0010","0010","0100","1010","1010","0111","0010","0010","0001","0010","0010","0011","0011","0100","0100","0100","0100","0100","0011","0100","0100","0100","0010","0001","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0100","0100","0100","0011","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0011","0101","1001","1001","1001","1001","0101","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0001","0010","0001","0010","0011","1000","0100","0011","0011","0011","0011","0011","0100","1000","0111","0110","0101","0101","0101","0101","0110","0111","0111","0111","0110","0101","0010","0001","0001","0001","0100","1000","1000","1000","0111","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0111","0110","0010","0001","0001","0001","0010","0100","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0010","0010","0011","0011","0011","0010","0001","0000","0010","0100","0101","0101","0101","0101","0101","0100","0101","0101","0110","0110","0110","0110","0111","0110","0011","0001","0010","0001","0001","0011","0110","0110","0110","0110","0110","0101","0011","0011","0110","0110","0110","0111","0110","0110","0101","0011","0010","0101","0111","0110","0110","0110","0110","0110","0110","0101","0100","0101","0101","0101","0101","0110","0110","0110","0110","0101","0110","0100","0001","0001","0010","0101","0110","0101","0101","0100","0100","0100","0101","0101","0110","0110","0010","0001","0001","0001","0001","0010","0110","0110","0110","0110","0110","0101","0100","0101","0110","0111","0110","0111","0011","0001","0001","0001","0010","0011","0110","0110","0101","0110","0100","0011","0011","0100","0101","0101","0100","0001","0010","1000","1000","0110","1000","1000","0110","0101","0101","0100","0101","0101","0101","1000","1100","0111","0110","1010","0100","0010","0111","0111","0111","0100","0011","0010","0100","0010","0001","0001","0000","0001","0011","0101","0111","1001","1000","1000","0111","0010","0001","0001","0001","0010","0010","0001","0001","0010","0100","0100","0100","0100","0011","0010","0011","0100","0101","1000","1000","0100","0011","0101","0101","0100","0010","0100","0101","0100","0101","0101","0100","0100","0100","0100","0100","0011","0011","0011","0100","0011","0101","0110","0100","0010","0011","0100","0011","0100","0100","0100","0011","0010","0011","0011","0011","0011","0010","0010","0011","0100","0101","0100","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0101","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0110","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0110","0110","0110","0101","0101","0101","0100","0100","0100","0100","0101","0110","0110","0110","0110","0110","0110","0110","0100","0100","0100","0101","0101","0100"),
("0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0110","0010","0011","0101","0101","0101","0100","0100","0100","0101","0100","0100","0101","0011","0110","0110","0101","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0110","0110","0111","0111","0110","0110","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0101","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0101","0011","0010","0010","0010","0010","0010","0011","0111","1000","1000","0011","0010","0011","0100","0101","1000","0111","0011","0001","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0001","0010","0010","0010","0011","0100","0100","0011","0011","0011","0011","0100","0101","0101","0101","0101","0110","0111","1001","1001","1001","1001","1000","0011","0010","0010","0010","0011","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0010","0010","0001","0101","1010","0110","0011","0011","0011","0011","0011","0100","1000","1000","0110","0101","0101","0101","0101","0110","0111","0111","0111","0110","0101","0010","0001","0001","0001","0100","1000","1000","1000","0111","0110","0110","0110","0101","0101","0101","0110","0110","0111","0111","0110","0110","0110","0010","0001","0001","0001","0010","0100","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0010","0010","0011","0011","0010","0010","0010","0001","0001","0011","0101","0101","0110","0101","0101","0100","0100","0101","0110","0110","0110","0110","0111","0101","0010","0001","0010","0010","0001","0010","0110","0110","0110","0101","0101","0101","0011","0011","0101","0110","0110","0111","0111","0101","0010","0001","0001","0001","0101","0110","0110","0110","0110","0111","0110","0101","0101","0110","0110","0110","0100","0101","0101","0110","0110","0110","0110","0010","0000","0001","0001","0011","0110","0110","0110","0101","0011","0011","0011","0100","0100","0101","0001","0001","0001","0001","0010","0010","0110","0110","0110","0110","0110","0101","0100","0100","0101","0110","0110","0110","0100","0001","0001","0010","0011","0101","0101","0110","0101","0101","0100","0011","0100","0100","0101","0101","0011","0001","0101","1001","0111","0111","0111","0101","0101","0110","0111","0111","0110","0110","0101","0110","1010","1011","0101","1001","1000","0010","0010","0111","0111","1000","0101","0011","0011","0001","0001","0001","0001","0001","0001","0001","0100","0111","0100","0100","0011","0010","0001","0001","0001","0011","0011","0001","0001","0010","0100","0100","0100","0100","0100","0100","0011","0010","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0100","0110","1000","0111","0111","0110","0100","0100","0100","0100","0100","0100","0110","0111","0111","0111","0110","0101","0110","0101","0100","0100","0101","0101","0101","0100","0101","0110","0110","0110","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0101","0100"),
("0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0010","0100","0100","0011","0100","0101","0101","0010","0010","0110","0101","0011","0011","0100","0110","1000","1000","0111","0010","0010","0010","0010","0100","0011","0010","0010","0001","0001","0010","0010","0010","0001","0010","0001","0001","0001","0001","0010","0010","0010","0010","0001","0001","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0101","0110","0110","0111","0101","0101","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0100","0110","1000","0111","0011","0010","0011","0010","0010","0011","0011","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0101","0100","0100","0101","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0011","0100","0110","0011","0010","0011","0010","0111","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","0110","0010","0010","0010","0010","0011","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","1000","1001","1000","0101","0011","0011","0011","0011","0101","0111","1000","0111","0101","0101","0101","0100","0110","0111","0110","0111","0110","0101","0010","0001","0001","0001","0011","0111","0111","1000","0110","0110","0110","0110","0101","0101","0101","0110","0110","0111","0111","0110","0111","0110","0010","0001","0001","0001","0010","0011","0100","0101","0110","0101","0101","0101","0101","0110","0110","0110","0111","0110","0011","0001","0011","0100","0010","0010","0001","0010","0001","0010","0101","0101","0110","0101","0110","0110","0101","0110","0110","0110","0111","0111","0111","0110","0010","0010","0001","0010","0010","0001","0101","0110","0110","0110","0100","0100","0011","0100","0110","0110","0111","1000","0111","0100","0010","0001","0001","0001","0011","0111","0111","0111","0110","0110","0100","0100","0100","0101","0101","0100","0011","0011","0100","0101","0101","0110","0101","0001","0001","0001","0010","0100","0111","0111","0111","0110","0011","0011","0011","0100","0100","0101","0001","0001","0001","0001","0010","0011","0110","0110","0110","0111","0110","0101","0100","0100","0100","0101","0101","0110","0100","0001","0001","0010","0100","0101","0110","0110","0110","0110","0100","0011","0100","0101","0110","0110","0011","0010","1000","1001","0110","1000","1000","0100","0100","0100","0110","0011","0101","0100","0101","0100","0111","1011","1000","0111","1010","0101","0001","0010","0110","1000","1000","0111","0010","0010","0001","0001","0001","0001","0001","0001","0011","0101","0010","0010","0001","0001","0001","0001","0001","0010","0100","0001","0001","0010","0011","0011","0011","0100","0011","0010","0010","0010","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0101","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0100","0110","1000","1000","0111","1000","0011","0010","0001","0001","0010","0011","0111","0111","1000","0111","0110","0110","0111","0111","0100","0010","0010","0001","0011","0011","0111","1000","0110","0111","0110","0111","0111","0100","0011","0010","0010","0011","0100","0111","0111","0110","0111","0101","0111","0111","0100","0011","0011","0011","0011","0011","0110","0111","0110","0110","0111","0110","0110"),
("0100","0100","0100","0100","0100","0100","0010","0010","0010","0010","0010","0001","0001","0001","0001","0100","0110","0101","1000","0111","0010","0001","0010","1000","1000","0110","0110","0111","1001","1011","1010","1001","0111","0100","0010","0010","0100","0101","0011","0010","0010","0001","0010","0001","0010","0001","0001","0010","0010","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0101","0110","0110","0111","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0101","0100","0010","0011","0010","0010","0010","0011","0100","0011","0010","0001","0010","0010","0011","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0101","0100","0100","0100","0100","0011","0010","0011","0100","0100","0100","0100","0100","0101","0110","0101","0110","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0101","0101","0010","0010","0010","0010","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0011","0001","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0110","0011","0010","0010","0001","0100","1010","1001","1001","1001","0011","0011","0011","0011","1000","1001","1001","1000","0110","0110","0101","0101","0110","0110","0110","0111","0110","0101","0010","0001","0010","0001","0011","1000","1001","1000","0111","0110","0111","0111","0110","0110","0110","0111","1000","1000","1000","1000","1000","0111","0010","0001","0001","0001","0010","0100","0101","0110","0101","0100","0100","0011","0011","0100","0100","0100","0100","0100","0010","0001","0010","0011","0010","0001","0000","0010","0001","0010","0100","0101","0111","0101","0110","0110","0101","0110","0101","0110","0110","0111","0111","0101","0010","0010","0000","0010","0010","0000","0101","0110","0110","0110","0101","0101","0100","0100","0110","0101","0110","0111","0111","0011","0010","0001","0001","0001","0010","0110","0111","0111","0110","0101","0101","0100","0100","0101","0101","0100","0100","0100","0100","0100","0101","0110","0101","0001","0001","0001","0010","0101","0111","0111","0110","0101","0011","0011","0011","0100","0101","0101","0001","0001","0001","0001","0010","0100","0110","0110","0110","0110","0110","0101","0101","0101","0110","0111","0110","0111","0101","0001","0001","0011","0101","0101","0111","1000","0111","0110","0101","0011","0100","0101","0110","0101","0011","0110","1010","0111","0111","0111","0110","0100","0101","0011","0101","0011","0101","0011","0101","0100","0101","1001","1011","0111","1001","1010","0100","0010","0010","0111","1001","0111","0110","0010","0001","0010","0001","0001","0001","0000","0110","0100","0001","0001","0001","0001","0001","0001","0010","0011","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","0101","0101","0110","0101","0010","0001","0010","0010","0010","0010","0001","0001","0010","0010","0001","0001","0001","0100","0110","1000","1000","0111","1000","0100","0100","0011","0010","0100","0100","1000","1000","1000","0111","0110","0110","1000","1000","0100","0011","0011","0010","0010","0001","0011","0101","0110","0110","0110","1000","0111","0100","0010","0001","0000","0010","0011","0110","0111","0110","0110","0110","1000","0111","0100","0010","0010","0001","0011","0010","0110","1000","0110","0110","0111","0111","0110"),
("0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0001","0001","0001","0001","0010","0111","1001","1001","0111","0001","0001","0010","0110","1000","1000","1000","1000","1000","1001","1001","1001","1000","0111","0101","0010","0010","0011","0011","0010","0010","0010","0001","0010","0010","0010","0001","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0011","0010","0010","0010","0101","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0101","0101","0110","0111","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0100","0100","0011","0011","0011","0100","0011","0011","0100","0101","0011","0011","0010","0001","0010","0011","0100","0100","0011","0011","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0011","0100","0100","0100","0100","0100","0011","0100","0011","0101","0101","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0011","0011","0011","0011","0011","0010","0010","0011","0100","0010","0010","0011","0011","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","0111","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1000","1000","0010","0010","0010","0010","0111","1010","1001","1000","1011","0101","0011","0011","0011","0100","0101","0101","0100","0011","0011","0011","0011","0101","0110","0110","0111","0110","0101","0010","0001","0001","0001","0011","1000","1000","1000","0111","0111","0110","0110","0101","0110","0101","0101","0110","0111","0111","0111","0110","0110","0011","0001","0001","0001","0010","0100","0101","0101","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0001","0001","0010","0011","0011","0010","0001","0010","0010","0010","0100","0101","0110","0110","0110","0101","0101","0101","0110","0110","0110","0110","0110","0100","0010","0010","0010","0010","0010","0010","0100","0110","0110","0110","0101","0101","0011","0100","0110","0110","0111","0111","0111","0101","0010","0010","0001","0010","0010","0101","0111","0111","0110","0110","0101","0101","0100","0100","0101","0100","0100","0100","0100","0101","0101","0101","0101","0001","0001","0010","0010","0101","0111","0111","0111","0101","0100","0011","0100","0101","0110","0101","0001","0001","0001","0010","0011","0100","0110","0111","0110","0110","0110","0101","0100","0101","0110","0110","0101","0111","0101","0001","0001","0011","0100","0101","0111","0111","0111","0111","0101","0011","0100","0100","0101","0101","0101","1010","1000","0101","1000","0100","0101","0101","0101","0010","0101","0100","0101","0011","0110","0101","0101","0101","1011","1001","0100","1010","0111","0010","0100","0011","0110","0111","0111","0111","0010","0010","0010","0001","0001","0010","1000","0011","0011","0100","0100","0010","0001","0001","0010","0010","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0101","0100","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","0110","1000","1000","0111","1000","0101","0100","0100","0100","0100","0101","1000","0111","0111","0111","0110","0110","1000","1000","0101","0100","0100","0100","0010","0000","0000","0011","0110","0110","0110","1000","1000","0101","0101","0011","0010","0100","0100","0010","0010","0010","0101","0110","1000","1000","0100","0011","0100","0011","0100","0100","0111","1000","0110","0110","0111","0110","0110"),
("0100","0100","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0011","0101","0101","0011","0001","0001","0010","0011","0011","0011","0100","0100","0101","0101","0101","0100","0100","0100","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0001","0001","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0100","0010","0011","0100","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0011","0110","0110","0110","0111","0111","0110","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0001","0011","0110","0101","0101","0011","0011","0011","0011","0011","0011","0101","0110","0011","0011","0011","0010","0010","0010","0010","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0011","0011","0011","0100","0100","0100","0011","0011","0100","0100","0011","0010","0011","0011","0111","1001","1001","1001","1001","1001","1001","1001","1000","1001","0100","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","1001","1010","1001","1001","1011","1001","0011","0011","0011","0011","0101","0111","0101","0100","0100","0011","0100","0101","0110","0110","0110","0110","0100","0010","0010","0010","0010","0100","0110","0101","0110","0101","0100","0100","0100","0100","0101","0100","0101","0110","0110","0110","0101","0101","0101","0011","0001","0001","0001","0010","0100","0101","0110","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0010","0001","0010","0011","0011","0010","0001","0001","0010","0010","0100","0101","0111","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0101","0011","0010","0010","0010","0010","0010","0100","0110","0110","0110","0110","0101","0011","0011","0101","0110","0111","0111","0110","0100","0011","0010","0001","0001","0001","0100","0110","0111","0110","0110","0110","0101","0100","0100","0101","0100","0100","0101","0101","0110","0101","0101","0110","0001","0001","0010","0011","0100","0110","0110","0101","0100","0011","0100","0100","0101","0110","0110","0001","0001","0001","0010","0100","0100","0110","0111","0110","0110","0110","0110","0101","0101","0110","0110","0110","0111","0101","0001","0001","0011","0101","0101","0111","0111","0111","0111","0101","0011","0100","0100","0101","0101","1000","1001","0110","0110","0110","0011","0110","0101","0011","0001","0100","0101","0101","0010","0101","0110","0101","0011","0111","1011","0110","0111","1011","0101","0011","0011","0001","0101","0111","1000","0111","0010","0001","0001","0000","0101","0111","0011","0100","0110","0101","0010","0001","0001","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0100","0100","0101","0100","0100","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0101","0110","0110","0100","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0011","0110","1000","1000","1000","1001","0101","0011","0010","0010","0010","0100","1000","1000","1000","0111","0110","0111","1000","1000","0101","0011","0011","0010","0001","0001","0001","0011","0111","0111","0110","0111","0110","0100","0100","0011","0010","0100","0100","0011","0011","0011","0100","0101","0111","0111","0100","0011","0011","0010","0011","0011","0110","1000","0110","0110","0111","0110","0110"),
("0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0011","0011","0010","0011","0011","0010","0100","0100","0100","0011","0010","0010","0011","0100","0011","0011","0100","0100","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0011","0010","0001","0001","0001","0001","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0110","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0011","0101","0101","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0110","0101","0011","0010","0001","0100","0110","0110","0110","0011","0100","0101","0100","0100","0100","1001","1000","0110","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0101","0101","0100","0101","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0111","1001","1000","1001","1001","1001","1001","1001","1000","0111","0010","0001","0010","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0100","0100","0010","0010","0010","0010","0110","1010","1010","1010","1001","1011","1011","0100","0011","0100","0100","0111","0111","0110","0101","0100","0100","0100","0101","0110","0111","0111","0110","0100","0010","0001","0010","0010","0011","0111","1000","1000","0110","0101","0101","0101","0101","0110","0110","0110","0111","0111","0111","0110","0110","0110","0011","0001","0001","0001","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0010","0001","0010","0100","0011","0010","0001","0001","0001","0001","0100","0101","0110","0101","0101","0100","0100","0101","0110","0110","0110","0110","0110","0100","0011","0010","0001","0001","0001","0001","0011","0101","0101","0101","0101","0101","0011","0011","0101","0110","0111","0111","0110","0100","0010","0010","0010","0001","0001","0100","0101","0110","0110","0110","0110","0101","0100","0100","0101","0100","0101","0101","0101","0110","0110","0111","0110","0001","0001","0010","0011","0100","0110","0110","0110","0101","0011","0100","0100","0101","0110","0110","0001","0001","0001","0010","0011","0101","0110","1000","1000","0111","0111","0110","0101","0100","0101","0101","0110","0111","0100","0001","0001","0011","0101","0101","0111","0111","0111","0111","0101","0011","0100","0100","0101","0101","0111","0111","0111","1000","0011","0100","0100","0101","0011","0010","0101","0101","0101","0001","0011","0110","0101","0100","0011","1010","1010","0101","1010","1001","0100","0010","0010","0010","0100","1001","0111","0111","0011","0001","0010","0111","0011","0101","0100","0011","0010","0001","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0100","0100","0110","0110","0110","0101","0101","0101","0101","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0001","0001","0001","0011","0101","0101","0100","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0111","0111","0110","0111","0101","0011","0100","0011","0100","0100","0101","0101","0101","0101","0100","0100","0101","0101","0100","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0110","0111","1000","0111","0111","0110","0111","0110","0110","0110","0111","0111","0111","0100","0011","0011","0011"),
("0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0001","0001","0001","0001","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0001","0001","0010","0010","0010","0100","0100","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0010","0010","0010","0010","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0011","0110","0110","0110","0101","0011","0100","0011","0011","0011","0011","0011","0101","0011","0010","0010","0010","0001","0001","0010","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0010","0100","1000","0110","0011","0011","0001","0101","1000","0110","0110","0011","0100","0110","0100","0010","0100","1010","1011","1010","1000","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","1000","1010","0101","0011","0010","0010","0100","0100","0101","0101","0011","0011","0100","0101","0100","0100","0101","0011","0011","0011","0011","0110","1001","1001","1001","1000","1000","1000","1000","1000","0100","0010","0011","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0011","0010","0010","0010","0010","0010","1000","1010","1010","1010","1001","1011","1100","1001","0100","0100","0110","0111","0111","0110","0101","0101","0100","0011","0101","0110","0111","0111","0110","0101","0010","0001","0001","0001","0011","1000","1001","1000","0111","0111","0110","0110","0101","0110","0110","0110","0111","0111","0111","0110","0110","0110","0011","0001","0001","0001","0010","0010","0010","0010","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0010","0001","0010","0011","0011","0010","0001","0001","0001","0001","0100","0100","0101","0101","0101","0100","0100","0101","0110","0110","0110","0110","0110","0101","0011","0010","0001","0010","0001","0001","0011","0110","0110","0110","0110","0101","0011","0011","0100","0111","0111","0111","0111","0100","0011","0010","0010","0001","0001","0100","0111","0111","0110","0110","0110","0101","0100","0100","0101","0101","0101","0101","0101","0101","0110","0111","0110","0001","0001","0010","0100","0101","0111","0111","0110","0101","0100","0100","0101","0101","0110","0110","0010","0001","0001","0010","0011","0100","0110","0111","1000","0111","0111","0110","0101","0101","0101","0101","0110","0111","0101","0001","0010","0011","0101","0101","0111","0111","0111","0111","0101","0100","0100","0101","0101","0101","0110","0110","1000","0111","0010","0101","0100","0110","0010","0010","0101","0011","0101","0010","0011","0110","0100","0110","0001","0110","1011","1000","1000","1011","0101","0001","0001","0001","0001","0100","0110","0011","0110","0011","0101","0110","0100","0110","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0011","0100","0110","0110","0110","0101","0100","0100","0011","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0001","0010","0001","0010","0001","0010","0010","0001","0001","0001","0011","0100","0100","0011","0100","0101","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0011","0100","0101","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0011","0010","0011","0011"),
("0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0010","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0100","0110","0101","0100","0100","0011","0011","0011","0011","0100","0011","0011","0011","0100","0100","0011","0010","0010","0100","0111","0110","0011","0010","0010","0010","0011","0101","0110","0110","0110","0110","0110","0110","0101","0011","0011","0011","0010","0100","0110","0100","0011","0011","0010","0100","0110","0101","0110","0011","0101","0101","0011","0010","0100","1010","1011","1011","1011","1010","0111","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0011","0011","0100","0100","0101","0100","0100","0100","0100","0011","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","1001","1011","1011","1011","0110","0011","0010","0011","0100","0101","0101","0101","0011","0100","0100","0100","0011","0100","0101","0011","0010","0010","0011","0110","1001","1000","1001","1000","1000","1000","1000","0111","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0001","0010","0010","0010","0100","1001","1010","1010","1010","0111","0101","0110","0110","0100","0011","0011","0100","0110","0101","0100","0100","1001","0111","1010","1010","1010","1001","0101","0100","0010","0010","0010","0010","0011","0101","0101","0101","0100","0100","0100","0011","0011","0111","0011","0011","0110","0111","0110","0110","0110","0111","0011","0001","0001","0001","0001","0001","0010","0011","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0010","0001","0010","0011","0011","0001","0001","0001","0001","0001","0100","0100","0101","0110","0101","0100","0100","0100","0101","0110","0110","0110","0110","0101","0011","0010","0001","0010","0001","0001","0100","0110","0110","0110","0101","0101","0011","0011","0101","0111","0111","0111","0110","0101","0100","0010","0010","0001","0001","0100","0111","0111","0110","0110","0110","0101","0100","0101","0101","0101","0101","0101","0101","0101","0110","0111","0110","0001","0001","0010","0100","0101","0110","0110","0110","0101","0100","0100","0101","0101","0101","0101","0010","0001","0001","0010","0100","0100","0110","0111","1000","1000","0111","0110","0101","0101","0101","0101","0101","0111","0101","0001","0010","0011","0101","0101","0111","0111","0111","0111","0101","0100","0101","0101","0110","0100","0100","0110","1000","0100","0100","0101","0101","0100","0001","0010","0101","0011","0110","0011","0010","0011","0100","0110","0011","0011","1001","1011","0101","1000","1001","0010","0001","0001","0010","0001","0100","0110","0011","0110","1000","0010","0111","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0100","0110","0110","0110","0110","0110","0110","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0010","0100","0101","0101","0101","0110","0110","0101","0110","1000","1000","0110","0100","0111","0111","0111","0100","0101","0101","0101","0100","0110","0110","0110","0110","0101","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0100","0100","0100","0110","0111","0111","0111","1000","1000","1000","1000","1000","1000","0111","1000","1000","0100","0011","0011","0011"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0010","0010","0011","0010","0010","0010","0001","0010","0010","0001","0001","0001","0010","0010","0010","0010","0100","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0101","0101","0101","0101","0100","0010","0001","0010","0010","0010","0011","0011","0011","0011","0101","0100","0011","0011","0100","0101","0010","0010","0100","0110","0110","0110","0100","0011","0100","0111","0110","0011","0011","0011","0011","0100","0101","0111","0111","0111","0110","0100","0110","0110","0101","0100","0011","0010","0011","0101","0110","0011","0011","0011","0100","0101","0011","0011","0100","0111","0011","0010","0011","0100","1001","1011","1011","1011","1011","1011","1001","0111","0101","0100","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0111","1001","1011","1011","1011","1011","1011","0110","0100","0100","0100","0101","0100","0101","0101","0100","0100","0100","0100","0011","0100","0101","0011","0010","0010","0011","0111","0101","0100","0100","0110","1000","1000","1000","0110","0001","0001","0001","0010","0011","0010","0010","0100","0110","0101","0101","0011","0010","0010","0010","0100","1001","1001","1000","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","1000","1010","1010","1001","0111","0101","0100","0010","0001","0010","0100","0011","0011","0011","0010","0010","0100","0110","0100","0110","1011","1100","0111","0010","0010","0010","0010","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0110","0110","0010","0010","0110","0111","0111","0110","0110","0110","0011","0001","0001","0010","0010","0011","0011","0011","0101","0110","0101","0101","0100","0101","0101","0101","0101","0101","0010","0001","0010","0100","0011","0011","0010","0011","0011","0001","0100","0100","0111","0110","0101","0100","0100","0100","0101","0111","0110","0101","0110","0101","0011","0010","0001","0001","0001","0001","0100","0110","0110","0110","0110","0101","0100","0011","0101","0111","1000","1000","0111","0101","0100","0011","0010","0001","0001","0100","0101","0110","0101","0101","0110","0101","0100","0110","0110","0101","0101","0110","0101","0101","0101","0111","0110","0001","0001","0010","0011","0100","0110","0110","0110","0101","0100","0100","0100","0100","0100","0101","0001","0001","0001","0010","0100","0100","0110","1000","0111","0110","0110","0101","0101","0101","0101","0100","0100","0111","0101","0001","0010","0011","0101","0101","0111","0111","0111","0111","0101","0100","0101","0101","0110","0100","0101","1001","0101","0100","0101","0110","0110","0011","0001","0001","0101","0100","0101","0010","0010","0100","0101","0110","0101","0011","0110","1011","1000","0100","1010","0110","0001","0010","0010","0010","0001","0011","0111","1000","1010","1000","1000","0010","0011","0011","0101","0100","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0001","0101","0110","0110","0110","0110","0110","0101","0011","0001","0010","0010","0001","0010","0011","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0011","0110","0110","0110","0110","0110","0110","0101","1010","1100","1100","0111","0111","1011","1100","1001","0101","1010","1100","1010","0101","0110","0110","0110","0110","0101","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0101","0111","0110","0110","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0100","0011","0011","0011"),
("0001","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0001","0010","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0101","0101","0011","0001","0001","0011","0101","0110","0111","0111","0110","0110","0101","0011","0010","0010","0011","0100","0100","0101","0101","0110","0100","0010","0100","0110","0101","0101","0100","0011","0011","0101","0110","0011","0011","0010","0100","0011","0010","0010","0110","0101","0100","0100","0100","0100","1010","1011","1011","1011","1011","1011","1011","1011","1001","0110","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0111","1010","1011","1011","1011","1011","1011","1011","1011","0101","0011","0100","0100","0100","0011","0100","0101","0100","0100","0100","0100","0100","0101","0101","0100","0010","0011","0011","0111","0100","0000","0001","0100","0101","0111","1000","0011","0001","0010","0001","0010","0010","0010","0001","1000","1011","1011","1011","0101","0010","0010","0010","0101","1010","1010","1010","1000","0010","0010","0010","0010","0010","0010","0001","0001","0010","0011","0011","0101","0101","0100","0110","1000","1000","1010","1010","1010","0101","0100","0101","0101","0001","0010","0011","0010","0011","0011","0010","0100","1001","0100","0000","0100","1010","1001","0100","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0010","0010","0010","0010","0110","0010","0001","0010","0011","0011","0011","0011","0011","0011","0010","0001","0001","0010","0011","0011","0011","0010","0011","0100","0100","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0011","0101","0100","0001","0100","0101","0111","0111","0110","0101","0101","0101","0110","0110","0110","0110","0110","0101","0100","0010","0001","0001","0001","0001","0100","0110","0110","0111","0110","0110","0101","0011","0100","0110","0111","0111","0111","0101","0011","0010","0001","0001","0001","0011","0110","0110","0101","0101","0110","0101","0100","0101","0101","0100","0100","0110","0101","0100","0100","0110","0110","0001","0001","0010","0011","0100","0110","0110","0110","0101","0100","0100","0101","0100","0101","0101","0011","0100","0100","0011","0011","0100","0110","1000","0110","0110","0110","0101","0100","0101","0101","0100","0100","0111","0110","0011","0011","0100","0101","0101","0110","0111","0110","0111","0101","0100","0110","0110","0110","0101","0101","0111","0010","0010","0101","0101","0111","0101","0100","0100","0101","0101","0101","0011","0011","0100","0111","0111","0101","0010","0010","1000","1011","0110","0111","1010","0011","0010","0010","0010","0001","0001","0100","1000","0110","1000","1000","0111","0110","0101","0100","0010","0100","0100","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0100","0100","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0110","0110","0110","0110","0110","0110","0101","0010","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0001","0010","0010","0010","0001","0010","0010","0010","0001","0010","0001","0001","0001","0010","0100","0110","0110","0110","0110","0110","0110","0110","1011","1100","1011","0110","1010","1011","1100","0111","1001","1100","1100","1010","0101","0110","0110","0110","0110","0100","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0000","0100","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","1000","0111","0111","0111","0111","0110","0011","0011","0011","0011"),
("0001","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0001","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0101","0011","0010","0011","0101","0100","0010","0010","0011","0100","0110","0111","0101","0101","0100","0110","0101","0110","0110","0110","0110","0100","0011","0101","0111","1000","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0101","0100","0011","0100","0100","0101","0100","0100","0101","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1001","0111","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0101","1000","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","0110","0100","0100","0100","0100","0011","0011","0100","0100","0101","0101","0100","0100","0101","0101","0100","0010","0011","0011","0111","0100","0001","0010","0001","0010","0110","0101","0010","0011","0010","0010","0010","0010","0010","0001","0111","1011","1010","1011","0101","0010","0010","0001","0101","1011","1011","1011","1000","0010","0011","0011","0100","0100","0011","0010","0010","0111","1010","1001","1010","1010","1001","1001","1001","0111","1011","1000","0100","0101","0101","0101","0101","0010","0010","0011","0011","0011","0011","0010","1000","1010","0101","0000","0101","1010","0110","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0100","0100","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0101","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0100","0010","0100","0101","0101","0101","0100","0100","0100","0100","0110","0111","0111","0110","0110","0101","0100","0010","0001","0001","0001","0001","0011","0110","0110","0101","0100","0100","0100","0011","0101","0110","0110","0111","0110","0101","0100","0010","0010","0001","0001","0100","0110","0111","0110","0110","0110","0110","0100","0100","0101","0100","0100","0110","0101","0101","0101","0110","0101","0001","0001","0010","0011","0100","0110","0111","0111","0110","0100","0011","0100","0100","0100","0100","0110","0110","1000","1000","0101","0100","0101","0110","0110","0111","0110","0110","0101","0101","0110","0101","0101","0111","0111","0111","0111","0110","0101","0101","0110","0110","0110","0110","0101","0010","0011","0011","0100","0100","0101","0011","0001","0010","0011","0011","0101","0011","0011","0100","0111","0111","0110","0011","0011","0011","0111","0100","0110","0010","0001","0100","1010","1001","0110","1010","1000","0010","0010","0011","0011","0011","0110","0100","0110","0111","0111","0111","0110","0100","0101","0101","0110","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0101","0101","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0101","0100","0001","0001","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0101","0110","0110","0110","0110","0110","0101","0101","1000","1000","0111","0100","1000","1001","1001","0101","1000","1001","1001","0110","0101","0110","0110","0110","0101","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0100","1000","1000","0111","0111","1000","1000","0111","1000","1000","0111","1000","1000","0111","0111","0111","0111","0110","0110","0101","0100","0101","0101"),
("0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0011","0010","0011","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0100","0101","0101","0011","0010","0011","0101","0011","0010","0011","0101","0111","1000","0111","1000","1001","1000","1001","1001","1001","1000","1011","1010","1000","1000","1010","1011","1011","1100","1011","1001","1000","1010","1010","1011","1010","1010","1011","0111","0101","0011","0100","0101","0101","0101","0100","0101","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","0111","0101","0100","0100","0101","0100","0101","0101","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0011","0011","0010","0010","0001","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0101","1000","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","0110","0100","0101","0110","0101","0001","0001","0010","0100","0101","0101","0101","0101","0101","0101","0100","0011","0010","0010","0100","0011","0001","0010","0010","0001","0001","0001","0010","0011","0010","0001","0010","0010","0010","0001","0111","1011","1011","1011","0101","0011","0011","0100","0101","1011","1100","1011","1010","1010","1011","1010","1001","1000","0110","0011","0010","0111","1000","1000","1000","0111","0111","0111","0110","0101","0110","0100","0011","0011","0010","0010","0010","0001","0010","0010","0010","0011","0010","0010","0011","0011","0010","0001","0011","0101","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0101","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0010","0010","0010","0100","0100","0100","0100","0100","0110","0110","0101","0101","0100","0100","0101","0110","0110","0110","0110","0101","0100","0010","0001","0001","0001","0001","0011","0110","0110","0101","0101","0101","0011","0010","0100","0110","0110","0111","0110","0101","0100","0011","0010","0001","0001","0100","0110","0110","0110","0110","0101","0101","0100","0100","0101","0100","0100","0100","0100","0101","0101","0110","0101","0001","0001","0011","0100","0100","0110","0111","0110","0101","0011","0010","0011","0011","0011","0100","0100","0101","1000","1001","1001","1000","0110","0111","0111","0111","0111","0110","0011","0011","0100","0100","0101","0110","1000","1000","1000","1000","0110","0101","0110","0110","0110","0110","0101","0011","0100","0100","0110","0101","0101","0011","0001","0011","0100","0101","0100","0010","0001","0001","0101","0011","0101","0001","0010","0010","0110","0100","0110","0011","0010","0010","0111","1011","1000","0110","1011","0101","0011","0100","0100","0111","0101","0010","1001","1011","1011","1011","1010","1010","1001","1000","1000","1000","0111","0110","0111","0110","0110","0111","0110","0110","0111","0110","0111","0111","0111","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0010","0001","0001","0001","0001","0011","0011","0010","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0010","0011","0110","0110","0110","0110","0110","0110","0101","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0100","0110","0110","0110","0110","0101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111"),
("0010","0010","0010","0010","0011","0010","0010","0011","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0011","0011","0011","0011","0011","0011","0100","0100","0101","0110","0100","0100","0011","0011","0100","0101","0111","1000","1001","1010","1001","1001","1001","0111","0111","0110","0110","0111","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1010","1001","1011","1010","0110","0101","0100","0100","0100","0100","0100","0100","0101","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1000","0101","0100","0101","0101","0101","0101","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0110","0111","1000","1000","1000","1000","1000","1000","1000","1000","0101","0110","1000","1000","1000","1000","1000","1000","1000","1000","1000","0110","0100","0011","0110","1001","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","0111","0101","0110","0110","0101","0010","0001","0011","0101","0101","0100","0100","0100","0011","0011","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0001","0001","0001","0001","0010","0010","0011","0011","0011","0001","0110","1011","1011","1011","1000","1001","1010","1011","0111","1011","1011","1011","1011","1010","1001","1000","0111","0110","0100","0001","0010","0100","0101","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0011","0100","0010","0001","0001","0010","0010","0010","0011","0011","0010","0010","0010","0010","0001","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0101","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0100","0100","0010","0010","0100","0100","0010","0100","0101","0110","0110","0101","0100","0100","0101","0101","0110","0110","0110","0101","0101","0100","0101","0101","0101","0110","0110","0101","0101","0101","0101","0110","0101","0011","0010","0100","0110","0110","0111","0111","0101","0100","0010","0010","0001","0001","0100","0101","0101","0101","0101","0100","0100","0011","0100","0101","0100","0100","0011","0011","0011","0100","0101","0110","0010","0010","0011","0100","0100","0110","0111","0110","0101","0011","0011","0011","0011","0100","0100","0100","0100","0111","0111","0111","0111","0110","0111","0111","0110","0110","0110","0100","0100","0101","0101","0110","0110","0101","0100","0100","0100","0100","0101","0111","0111","0110","0110","0100","0011","0100","0101","0110","0101","0101","0011","0001","0100","0101","0101","0011","0010","0010","0010","0101","0011","0101","0010","0010","0010","0101","0101","0110","0100","0001","0001","0011","1010","1001","0010","1000","1001","0110","0110","0111","1000","0011","0011","1001","1100","1011","1100","1100","1100","1011","1011","1010","1001","1000","0101","0111","0110","0110","1000","1000","1000","1000","0111","1001","1000","1000","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0001","0001","0001","0010","0011","0100","0011","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0011","0010","0001","0001","0001","0010","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0011","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0011","0010","0010","0010","0011","0011","0011","0100","0100","0100","0011","0100","0100","0011","0011","0011","0010","0011","0011","0011"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0100","0101","0110","0101","0101","0111","0111","1000","1000","1001","1001","1001","1010","1010","1001","1001","1000","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1000","0110","0101","0101","0100","0011","0100","0100","0100","0100","0101","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","0111","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0011","0011","0010","0010","0011","0100","0101","0110","0111","1000","1000","1001","1001","1001","1001","1001","0110","0110","1001","1001","1001","1001","1001","1001","1001","1001","0110","0010","0101","1001","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","0111","0101","0101","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0101","0100","0100","0100","0011","0010","0010","0011","0010","0001","0001","0001","0011","0100","0100","0101","0100","0100","0011","0110","1010","1100","1010","1001","1001","0111","0100","1000","1011","1100","1001","0101","0101","0101","0101","0100","0011","0010","0010","0100","0100","0100","0100","0100","0100","0101","0100","0101","0100","0100","0010","0010","0011","0011","0010","0001","0001","0010","0010","0011","0011","0011","0011","0011","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0011","0100","0011","0100","0010","0100","0110","0101","0101","0101","0101","0101","0101","0110","0111","0110","0011","0011","0011","0011","0100","0111","0111","1000","0111","0101","0101","0101","0100","0101","0011","0010","0100","0101","0110","0111","0110","0101","0100","0011","0010","0001","0010","0100","0110","0101","0101","0101","0100","0100","0100","0101","0101","0100","0100","0100","0011","0100","0101","0101","0110","0101","0110","0100","0100","0100","0110","0110","0101","0100","0100","0100","0100","0100","0100","0101","0100","0100","0110","0111","0111","0111","0111","0111","0110","0101","0110","0101","0100","0100","0110","0101","0110","0110","0101","0100","0100","0100","0100","0101","0111","0111","0111","0111","0100","0011","0100","0101","0101","0101","0101","0011","0001","0101","0110","0101","0010","0010","0010","0010","0101","0100","0101","0010","0011","0010","0100","0101","0101","0101","0001","0001","0001","0110","1011","0111","0101","1010","0111","1001","1000","0101","0100","0011","0110","1000","1000","1001","1001","1001","1001","1010","1010","1010","1001","0100","0010","0010","0101","0111","1000","0111","1000","1000","1001","1000","0110","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0001","0001","0001","0010","0010","0011","0011","0010","0001","0010","0001","0001","0001","0001","0010","0001","0001","0001","0010","0001","0010","0011","0010","0001","0001","0001","0010","0101","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001"),
("0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0011","0011","0011","0100","0100","0100","0011","0101","0101","0110","0111","1000","1001","1001","1010","1001","1001","1010","1001","1001","1001","1001","1010","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1100","1001","0101","0100","0010","0010","0010","0100","0100","0100","0100","0101","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1001","0101","0110","0011","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0001","0000","0000","0000","0000","0011","0110","0110","0110","0110","0110","0110","0110","0100","0101","0111","0111","0111","0110","0110","0110","0110","0110","0110","0101","0111","1010","1001","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","0011","0010","0010","0001","0001","0001","0001","0010","0001","0010","0011","0100","0100","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0011","0101","0111","0110","0101","0101","0100","0100","0011","0110","1011","1000","0100","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0010","0010","0011","0010","0001","0001","0010","0010","0011","0011","0011","0011","0011","0010","0001","0001","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0100","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0101","0110","1000","1000","1000","0111","0111","0111","0110","0100","0011","0011","0011","0011","0011","0010","0011","0100","0101","0101","0101","0010","0100","0110","0101","0101","0101","0101","0110","0111","0110","0101","0011","0011","0011","0011","0100","0100","0100","0101","0101","0110","0110","0101","0100","0110","0100","0010","0100","0101","0110","0110","0110","0101","0100","0010","0011","0011","0011","0101","0110","0101","0101","0101","0101","0100","0100","0101","0101","0101","0100","0100","0100","0101","0101","0101","0110","1000","1000","0111","0110","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0110","0100","0100","0110","0111","0110","0111","0111","0111","0111","0101","0110","0110","0100","0100","0110","0101","0110","0110","0101","0101","0101","0101","0100","0101","0111","0111","0111","0110","0100","0011","0100","0101","0101","0101","0110","0100","0011","0110","0100","0100","0010","0010","0010","0001","0100","0100","0101","0010","0101","0011","0100","0111","0110","0111","0010","0010","0010","0011","1001","1001","0110","1000","1010","1000","0101","0101","0011","0011","0100","0110","0111","1010","1010","1010","1000","0101","0110","1010","1001","0101","0010","0011","0100","0101","0100","0011","0111","0111","0110","0101","0100","0100","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0010","0001","0010","0001","0001","0001","0010","0010","0001","0010","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0010","0011","0010","0001","0001","0001","0010","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001"),
("0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0101","0110","0111","1000","1000","1001","1001","1001","1010","1001","1000","1000","1001","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","0111","0101","0011","0010","0010","0011","0100","0100","0100","0100","0100","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1001","0100","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0001","0000","0000","0000","0000","0100","0110","0110","0110","0110","0111","0111","0111","0101","0101","0111","0111","0111","0111","0110","0110","0110","0110","0111","0111","0100","0100","0100","1001","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1011","1010","1010","1010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","0101","0100","0011","0010","0001","0001","0001","0010","0010","0010","0010","0010","0001","0010","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0010","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0011","0010","0010","0011","0011","0101","0010","0010","0010","0011","0011","0011","0010","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","1000","1000","1011","1011","1010","1010","1010","1001","0110","0100","0011","0011","0010","0011","0010","0011","0100","0101","0101","0110","0101","0110","0010","0100","0110","0100","0101","0110","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0110","0110","0101","0110","0111","0101","0100","0101","0101","0110","0110","0110","0101","0101","0101","0101","0111","0110","0101","0110","0101","0101","0101","0101","0100","0011","0100","0100","0011","0100","0100","0100","0110","0101","0110","0111","0111","0111","0111","0111","0110","0110","0110","0101","0100","0100","0100","0101","0101","0110","0111","0100","0010","0010","0101","0110","0111","1000","1000","0111","0111","0111","0110","0101","0101","0110","0101","0110","0111","0101","0100","0100","0011","0011","0101","0110","0110","0110","0110","0101","0011","0100","0100","0101","0100","0101","0100","0100","0100","0011","0011","0010","0010","0010","0010","0110","0110","0111","0011","0100","0011","0011","0110","0011","0101","0100","0010","0010","0010","0110","0110","0011","0011","0110","0100","0011","0011","0011","0100","0011","0101","0011","0100","0100","0100","0011","0011","0011","1001","1001","0011","0001","0011","0100","0011","0011","0011","0011","0011","0010","0011","0010","0011","0100","0100","0101","0101","0110","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0110","0011","0010","0010","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0010","0001","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0101","0011","0010","0011","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001"),
("0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0110","0100","0100","0101","0101","0110","0110","0110","0111","0111","0110","0110","0110","0110","0111","0110","0111","0110","0101","0101","0110","0101","0101","0101","0101","0101","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0101","0101","0111","0100","0100","0011","0011","0011","0100","0110","0110","0100","0101","1001","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1000","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0011","0010","0010","0001","0001","0001","0001","0100","0110","0110","1000","1000","1001","1000","1000","0101","0101","0111","0111","1000","1000","1000","1001","1000","1000","1000","0111","0111","0100","0011","1000","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","0101","0100","0100","0011","0011","0011","0010","0010","0011","0010","0010","0010","0100","0101","0100","0011","0011","0010","0011","0010","0011","0011","0010","0010","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0001","0010","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0100","0011","0010","0010","0011","0011","0011","0011","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0110","1011","1011","1011","1011","1001","1010","1010","1000","0100","0100","0100","0011","0011","0100","0010","0100","0101","0101","0110","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0110","0101","0011","0100","0100","0100","0011","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0110","1000","0110","0100","0101","0101","0110","0110","0101","0100","0100","0100","0101","0100","0101","0010","0001","0100","0101","0110","0101","0100","0100","0100","0100","0010","0100","0100","0101","0100","0100","0100","0100","0100","0110","0111","0011","0001","0001","0011","0110","0111","1000","1000","1000","0111","0111","0110","0101","0101","0101","0101","0101","0110","0100","0011","0010","0011","0011","0101","0110","0110","0110","0101","0100","0011","0100","0100","0100","0100","0110","1000","1000","1000","1000","0100","0011","0011","0011","0011","0110","0011","0110","0011","0010","0011","0100","0100","0011","0011","0100","0011","0011","0010","0100","0101","0011","0011","0010","0010","0010","0010","0011","0111","0111","1010","0110","0110","0100","0100","0011","0011","0011","1000","1000","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0100","0100","0100","0100","0100","0011","0100","0101","0101","0110","0110","0110","0110","0110","0101","0011","0010","0100","0101","0010","0010","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0010","0010","0100","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001"),
("0010","0011","0010","0010","0010","0010","0010","0011","0011","0100","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0110","0101","0100","0101","0101","0101","0110","0110","0110","0110","0101","0110","0111","0110","0111","0111","0111","0111","0110","0110","0111","0110","0110","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0111","0101","0011","0100","0100","0100","0101","0100","0100","0100","0100","0100","0110","1101","1001","0100","0100","1001","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1000","0011","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0010","0010","0100","0011","0011","0010","0001","0001","0001","0001","0100","0110","0110","1000","0011","0011","0011","1000","0110","0101","0111","1000","1001","0011","0011","0100","0011","0011","0111","1000","0111","0101","0100","1000","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","0101","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0011","0100","0101","0101","0101","0101","0100","0011","0010","0011","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0100","0011","0010","0010","0011","0011","0011","0011","0011","0111","0111","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0111","1000","1010","1011","1011","1010","1010","1010","0110","0011","0011","0011","0011","0100","0011","0011","0100","0101","0101","0110","0110","0110","0101","0110","0111","0100","0100","0110","0110","0110","0110","0110","0101","0100","0100","0100","0100","0100","0101","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0101","0101","0110","0110","0110","0101","0101","0100","0101","0101","0100","0100","0011","0001","0001","0010","0100","0011","0011","0101","0111","0110","0011","0001","0011","0100","0011","0010","0010","0100","0100","0110","0111","0010","0001","0001","0010","0101","0111","1000","1000","0111","0111","0111","0101","0101","0100","0101","0100","0101","0110","0101","0011","0011","0011","0100","0101","0110","0110","0110","0110","0101","0011","0100","0100","0100","0100","0111","1011","1100","1100","1011","0100","0010","0010","0011","0011","0100","0010","0101","0011","0010","0010","0010","0011","0100","0010","0101","0010","0010","0010","0011","0101","0011","0010","0010","0011","0010","0100","0101","0110","0111","1000","0110","0110","0101","0100","0101","0101","0100","0100","0011","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0001","0010","0010","0011","0100","0100","0100","0011","0011","0100","0011","0100","0101","0101","0110","0110","0110","0110","0101","0100","0101","0100","0001","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0001","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0010","0001","0001","0011","0011","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0101","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0010","0100","0011","0010","0100","0011","0001","0001","0001","0001","0001","0001"),
("0010","0010","0010","0010","0010","0010","0011","0011","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0101","0110","0110","0110","0100","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0101","0101","0101","0100","0111","0101","0110","0111","0101","0110","0110","0110","0110","0111","0101","0011","0100","0100","0100","0100","0101","0101","0100","0100","0100","0111","1000","0101","0101","0100","1001","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1001","0100","0101","0101","0110","0101","0101","0101","0101","0011","0011","0110","0011","0001","0100","0101","0110","0011","0010","0100","0011","0011","0010","0001","0001","0001","0001","0100","0110","0110","1000","0010","0001","0001","0111","0110","0101","0111","1000","1000","0010","0001","0001","0001","0000","0110","0111","0111","0101","0101","1000","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1011","1010","0101","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0010","0011","0011","0100","0011","0010","0011","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0100","0011","0010","0011","0011","0011","0011","0011","0010","0010","0010","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0101","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0011","0110","0100","0010","1000","1100","1011","1011","1011","1001","0101","0011","0011","0011","0011","0011","0011","0011","0101","0101","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0111","0110","0100","0110","0110","0110","0111","0111","0111","0111","0111","0111","1000","1000","1000","0110","0101","0110","0110","0110","0101","0101","0100","0101","0101","0010","0001","0001","0001","0001","0001","0001","0001","0010","0011","0101","0100","0010","0001","0010","0011","0000","0000","0010","0100","0100","0101","0110","0010","0001","0001","0010","0101","0110","0111","0111","0111","0110","0111","0101","0101","0100","0100","0100","0110","0110","0101","0011","0010","0011","0101","1000","1000","1000","1000","0111","0101","0011","0100","0100","0100","0100","0100","1010","1100","1100","1011","0101","0101","0101","0011","0011","0101","0100","0011","0011","0011","0011","0011","0011","0100","0011","0011","0010","0010","0011","0101","0101","0011","0010","0010","0011","0011","0100","0101","0101","0100","0101","0011","0011","0010","0010","0011","0100","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0010","0001","0001","0001","0010","0001","0010","0011","0100","0100","0011","0011","0011","0100","0100","0100","0100","0101","0110","0110","0101","0101","0101","0101","0011","0001","0010","0010","0010","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0010","0010","0010","0001","0010","0010","0010","0001","0001","0001","0001","0001","0011","0100","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0010","0011","0110","0110","0110","0110","0110","0101","0011","0011","0011","0011","0010","0010","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0100","0011","0011","0010","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0110","0111","0110","0111","0100","0001","0001","0001","0001","0011","0100"),
("0010","0010","0010","0010","0011","0010","0011","0100","0011","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0110","0110","0100","0101","0101","0110","0111","0111","0111","0111","0111","0110","0111","0111","0111","1000","0111","0110","0111","0111","0111","0110","0011","0011","0011","0101","1000","0110","1001","0111","0101","0101","0101","0100","0100","0111","0101","0011","0100","0100","0101","0101","0101","0101","0100","0100","0011","0011","0011","0010","0010","0001","0110","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1000","0100","0110","0110","0110","0110","0011","0011","0110","0001","0011","0110","0011","0001","0101","0110","0110","0010","0010","0100","0100","0011","0010","0001","0001","0001","0001","0100","0110","0110","1000","0010","0001","0001","0111","0110","0101","0111","0111","1001","0010","0001","0001","0001","0001","0110","0111","0111","0101","0100","1000","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","0101","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0010","0011","0011","0011","0010","0011","0011","0011","0001","0001","0001","0001","0001","0001","0010","0100","0011","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0011","0100","0100","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0100","0010","0001","0011","0100","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0011","1001","0101","0011","1000","1011","1010","1010","1010","0101","0100","0011","0010","0011","0011","0100","0100","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0100","0100","0110","0110","0110","0101","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0111","0110","0110","0110","0111","0101","0100","0110","0110","0110","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0101","0101","0110","0101","0101","0101","0100","0101","0101","0011","0001","0001","0001","0000","0001","0000","0000","0011","0011","0001","0010","0001","0001","0001","0001","0000","0001","0001","0010","0011","0101","0110","0011","0001","0001","0010","0011","0110","0111","0111","0111","0110","0110","0101","0101","0100","0100","0011","0101","0101","0100","0001","0001","0010","0110","1100","1100","1100","1010","0110","0101","0010","0011","0011","0100","0101","0101","1010","1100","1011","1011","0110","0110","0101","0100","0011","0011","0011","0010","0011","0010","0011","0011","0010","0011","0011","0011","0010","0010","0011","0010","0011","0011","0011","0010","0011","0100","0100","0101","0100","0010","0010","0010","0100","0100","0100","0100","0100","0010","0010","0010","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0101","0101","0101","0101","0100","0100","0011","0001","0010","0001","0001","0001","0001","0001","0001","0001","0011","0010","0001","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0001","0001","0011","0100","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0010","0010","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0010","0010","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0010","0011","0010","0010","0100","0010","0001","0001","0010","0010","0011","0011","0010","0010","0001","0010","0010","0001","0111","1000","1000","0111","0100","0001","0001","0001","0001","0101","0111"),
("0010","0010","0010","0010","0011","0101","0101","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","1000","0111","0111","1000","1000","1000","1001","0111","0011","0110","0111","0111","0111","0111","0011","0011","0100","0101","0101","0100","0100","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0011","0100","0100","0011","0011","0010","0010","0001","0010","0010","0010","0010","0001","0101","1001","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1001","0100","0110","0110","0110","0110","0010","0100","0110","0010","0011","0111","0100","0001","0101","0111","0110","0011","0010","0101","0100","0011","0010","0001","0001","0001","0001","0100","0110","0110","1000","0010","0001","0001","0111","0110","0101","0111","0111","1001","0010","0001","0001","0001","0001","0110","1000","0111","0101","0100","0111","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","0101","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0001","0001","0010","0010","0001","0011","0001","0001","0010","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0011","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0101","0011","0011","0100","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0001","0010","0010","0010","0011","0110","0111","0101","0100","0101","0111","0101","0100","0100","0100","0100","0100","0011","0100","0101","0101","0011","0100","0101","0110","0110","0110","0110","0110","0110","0111","0110","0100","0100","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0100","0101","0011","0011","0101","0101","0010","0100","0101","0100","0101","0101","0100","0010","0001","0001","0001","0000","0000","0001","0001","0010","0010","0001","0010","0010","0001","0000","0001","0001","0001","0001","0010","0110","0110","0011","0001","0001","0001","0010","0101","0111","0111","0111","0110","0110","0101","0011","0010","0011","0101","0101","0110","0100","0001","0010","0010","0110","1100","1100","1101","1010","0110","0101","0011","0100","0100","0101","0100","0101","1010","1011","1000","0111","0100","0100","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0011","0100","0101","0100","0010","0010","0010","0001","0001","0010","0101","0100","0100","0100","0010","0010","0010","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0011","0010","0011","0011","0010","0011","0011","0011","0101","0101","0101","0101","0100","0011","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0011","0100","0100","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0010","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0110","0101","0101","0010","0010","0010","0010","0001","0110","1000","1000","0101","0010","0001","0001","0001","0001","0110","0111"),
("0010","0011","0011","0100","0011","0100","0100","0100","0100","0100","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0101","0011","0011","0011","0100","0101","0111","0111","1000","1000","1000","1001","0110","0010","0011","0110","0111","0110","0110","0101","0011","0011","0101","0100","0011","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","1000","1001","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1001","0100","0111","0111","0111","0110","0011","0100","0110","0010","0011","0111","0100","0010","0101","0111","0110","0011","0010","0101","0100","0011","0010","0001","0001","0001","0001","0100","0110","0110","1000","0011","0001","0001","0111","0110","0101","0111","0111","1001","0011","0001","0001","0001","0001","0110","1000","0111","0101","0100","1000","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","0101","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0001","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0010","0011","0011","0100","0011","0010","0001","0010","0010","0001","0011","0010","0010","0001","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0011","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0100","0010","0011","0011","0010","0010","0010","0011","0011","0100","0100","0100","0011","0011","0100","0100","0101","0101","0110","0101","0100","0011","0100","0100","0100","0011","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0100","0101","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","1000","0111","0010","0001","0001","0001","0011","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0011","0001","0001","0001","0001","0001","0001","0011","0100","0010","0001","0001","0001","0001","0100","0101","0101","0110","0101","0101","0101","0011","0100","0100","0101","0110","0111","0101","0001","0010","0010","0110","1010","1001","1000","1000","0110","0100","0011","0100","0100","0101","0100","0100","0101","0100","0110","0101","0010","0010","0011","0010","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0011","0010","0001","0010","0010","0010","0001","0001","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0100","0100","0100","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0101","0101","0100","0100","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0011","0100","0100","0100","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0011","0010","0010","0010","0100","0100","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0001","0001","0001","0010","0010","0011","0011","0010","0001","0001","0001","0001","0001","0010","0010","0001","0010","1000","1000","0111","0110","0110","0110","0110","0110","0111","1000","1000","0110","0011","0100","0100","0011","0011","0110","1000"),
("0011","0011","0011","0011","0010","0011","0100","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0101","0101","0101","0101","0101","0110","0100","0100","0011","0011","0110","1000","1000","1000","1001","1001","0110","0100","0011","0101","0110","0101","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","1000","1000","1001","1010","1010","1010","1010","1010","1011","1011","1011","1011","1001","0101","0111","0111","0111","0111","0011","0100","0111","0010","0100","0111","0100","0010","0110","0111","0111","0101","0011","0101","0100","0011","0010","0001","0001","0001","0001","0011","0110","0110","1000","0011","0001","0001","0111","0110","0101","0111","0111","1001","0010","0001","0001","0001","0001","0110","1000","0111","0101","0100","1000","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","1010","1011","1010","0101","0011","0100","0100","0100","0100","0011","0011","0011","0011","0010","0010","0001","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0001","0011","0010","0010","0010","0010","0001","0001","0001","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0100","0100","0010","0010","0011","0100","0100","0100","0100","0100","0100","0011","0011","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0100","0010","0010","0011","0011","0011","0011","0010","0001","0001","0001","0010","0010","0001","0001","0010","0011","0100","0011","0101","0100","0011","0100","0100","0011","0100","0100","0101","0101","0100","0100","0101","0110","0100","0100","0100","0011","0011","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0101","0011","0100","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0110","0110","0110","0111","0111","0111","0110","0111","0111","0111","1000","0111","0100","0011","0011","0011","0011","0011","0010","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0001","0001","0100","0101","0011","0001","0001","0001","0001","0011","0111","1000","1000","1001","1000","0101","0100","0100","0101","0101","0110","0111","0101","0001","0010","0010","0110","1010","1001","1001","1010","1000","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0010","0010","0010","0010","0010","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0010","0001","0010","0001","0001","0010","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0010","0100","0100","0011","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0101","0101","0101","0110","0110","0110","0110","0101","0001","0001","0010","0010","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0010","0010","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","1000"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0010","0011","0011","0011","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0010","0011","0101","0110","0101","0110","0110","0101","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0010","0010","0101","1000","1000","1000","1001","1010","0110","1001","1010","1010","1010","1011","1011","1001","0101","0111","0111","0111","0111","0011","0100","0111","0011","0100","0111","0100","0010","0110","0110","0110","0110","0100","0100","0011","0011","0011","0011","0100","0100","0010","0011","0110","0110","1000","0011","0000","0001","0111","0110","0101","0111","0111","1000","0100","0010","0001","0001","0001","0101","1000","0111","0101","0100","1000","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","0101","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0001","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0001","0010","0010","0010","0001","0001","0011","0011","0001","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0111","1000","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0101","0100","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0010","0011","0100","0101","0110","0110","0110","0101","0100","0011","0101","0111","1000","1000","1000","0111","1010","1010","1010","0101","0100","0110","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0101","0101","0101","0011","0011","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0101","0100","0011","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","0110","0100","0100","0101","0101","0101","0100","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0001","0010","0110","0111","0011","0010","0001","0001","0001","0010","0111","1101","1101","1100","1010","0101","0100","0101","0101","0101","0101","0111","0101","0010","0011","0011","0011","1001","1101","1100","1100","1001","0100","0111","0111","0110","0101","0100","0100","0011","0011","0011","0011","0010","0010","0011","0010","0010","0001","0001","0010","0010","0010","0001","0011","0011","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0010","0010","0010","0001","0010","0010","0010","0001","0010","0100","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0010","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0011","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0010","0110","1000","0011","0110","0110","0110","0110","0101","0010","0001","0001","0010","0001","0001","0001","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0011","1000","1000","0111","0110","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","1000"),
("0001","0010","0011","0011","0011","0010","0001","0001","0001","0001","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0001","0001","0010","0011","0100","0101","0101","0101","0101","0101","0100","0011","0011","0001","0000","0001","0001","0001","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0010","0010","0101","1000","1000","1000","1001","1001","0110","1001","1010","1010","1010","1010","1011","1001","0110","1000","1000","0111","0111","0011","0101","0111","0101","0100","0111","0100","0010","0101","0110","0010","0001","0010","0110","1000","1000","1001","1001","1001","1001","0111","0100","0101","0101","0110","0011","0010","0010","0110","0110","0100","0111","0111","1000","0111","0011","0001","0001","0000","0110","1000","0111","0101","0100","0111","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1011","0101","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0001","0010","0011","0010","0001","0001","0011","0011","0011","0010","0010","0101","0101","0101","0101","0101","0101","0101","0101","0111","0111","0110","0101","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0110","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0111","0110","0101","0101","0101","0011","0111","0011","0011","0011","0100","0100","0101","0011","0010","0100","0111","1001","1000","1010","0111","1011","1010","1011","0111","0110","0110","0101","0100","0100","0100","0100","0101","0101","0101","0110","0110","0101","0110","0101","0100","0011","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0101","0101","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0111","0111","0111","0111","1000","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0110","0100","0010","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0110","0111","0011","0001","0001","0001","0010","0101","0110","1010","1100","1011","1010","1001","1001","0111","0101","0101","0101","0101","0101","0101","0101","0100","0011","1001","1100","1100","1100","1001","0100","1000","1100","1011","0101","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0010","0101","0010","0010","0010","0010","0001","0010","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0011","0011","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0011","0100","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0101","0010","0110","1010","0101","0011","0100","0100","0100","0100","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0011","1000","1000","1000","0110","0110","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111"),
("0010","0010","0011","0110","0110","0101","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0011","0100","0100","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0101","0100","0100","0100","0100","0011","0001","0010","0011","0011","0100","0101","0101","0101","0101","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0101","0111","1000","1000","1001","1001","1001","1010","1010","1010","1010","1010","1000","0111","0110","0110","0101","0111","0110","0011","0010","0010","0010","0100","0111","0111","0110","1000","1000","0101","0010","0011","1000","1010","1010","1001","1001","1001","1001","1010","1001","0110","0101","0101","0101","0101","0101","0110","0101","0100","0111","0111","1001","0011","0001","0001","0001","0001","0101","1000","0111","0101","0100","0111","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","0101","0011","0011","0011","0011","0100","0100","0100","0011","0011","0010","0010","0001","0001","0001","0001","0011","0100","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0100","0100","0011","0010","0001","0010","0010","0001","0000","0001","0011","0011","0011","0010","0011","0101","0101","0111","0111","0100","0101","0101","0110","0111","0110","0101","0100","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","1000","0110","0110","0101","0101","0100","1001","0010","0001","0001","0010","0110","0111","0101","0101","0111","0111","0110","0111","1010","0111","1000","1010","1011","0111","0110","0110","0110","0101","0100","0100","0101","0101","0110","0110","0110","0110","0110","0101","0101","0100","0100","0100","0101","0110","0101","0101","0110","0110","0110","0110","0100","0001","0001","0001","0010","0101","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0111","0111","0101","0011","0010","0001","0001","0001","0101","0110","0110","0110","0101","0100","0011","0011","0010","0010","0001","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0010","0001","0001","0001","0011","1010","1011","1010","1000","1001","1100","1100","1100","1000","0100","0101","0100","0100","0101","0100","0101","0100","0100","1001","1100","1100","1100","1001","0100","1001","1100","1010","0100","0011","0011","0011","0010","0010","0010","0011","0010","0010","0011","0010","0010","0001","0001","0001","0001","0100","0110","0011","0010","0011","0010","0010","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0010","0001","0001","0010","0010","0001","0010","0010","0010","0001","0001","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0001","0010","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0010","0100","0110","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0110","1010","1001","1000","1001","1001","1001","0101","0010","0001","0001","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000"),
("0010","0010","0010","0100","0101","0100","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0101","0100","0001","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0100","0100","0011","0011","0011","0100","0011","0011","0011","0011","0010","0011","0100","0011","0011","0011","0010","0010","0010","0011","0011","0100","0100","0100","0101","0101","0101","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0101","0111","1000","1000","1001","1001","1001","1010","1010","1010","1010","1010","0101","0010","0010","0010","0011","0111","0111","0110","0100","0010","0001","0110","1010","1010","1010","1010","1001","1000","0111","0111","1000","1000","1001","1001","1001","1001","1001","1010","1010","1010","1000","0110","0101","0110","0110","0111","0101","0100","0111","0111","1001","0011","0001","0001","0001","0000","0101","1000","0110","0101","0011","0110","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","0110","0011","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0001","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0100","0100","0011","0010","0001","0010","0010","0001","0001","0010","0001","0010","0011","0010","0011","0100","0101","0101","0011","0011","0011","0100","0110","0111","0110","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","0110","0100","0100","0100","1001","0111","0111","0110","0110","1001","1100","1010","1010","1010","0011","0010","0011","0100","0100","0101","1000","1001","0110","0101","0011","0011","0100","0100","0100","0101","0110","0110","0110","0111","0110","0110","0110","0110","0011","0100","0011","0010","0011","0111","1000","1000","1000","0111","1000","0111","0110","0101","0101","0101","0111","0110","0111","0111","0110","0110","0111","0110","0110","0110","0110","0110","0111","0111","0111","0110","0001","0001","0001","0001","0001","0011","0101","0101","0100","0011","0010","0011","0011","0010","0010","0001","0001","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0101","1011","1100","1100","0101","1001","1101","1100","1100","1000","0100","0100","0101","0101","0101","0101","0101","0101","0100","1001","1100","1100","1100","1001","0100","1000","1010","0110","0100","0010","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0001","0001","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0010","0010","0011","0010","0010","0001","0010","0011","0011","0010","0010","0011","0010","0010","0011","0011","0010","0010","0011","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0001","0001","0010","0001","0010","0001","0001","0010","0010","0010","0001","0001","0010","0010","0010","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0101","1010","1000","1000","1001","1001","1001","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0100","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0010","0011","0011","0010","0001","0011","0010","0011","0100","0011","0011","0011","0101","0110","0110","0110","0011","0010","0010","0011","0010","0001","0001","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0101","0111","0111","1000","1000","1001","1001","1001","1010","1010","1010","1010","0110","0001","0010","0010","0100","1000","1001","1001","1000","0110","0101","0111","1001","1001","1001","1010","1001","1010","1001","1001","1001","1001","1000","1000","1001","1010","1010","1010","1010","1010","1010","1001","0111","0100","0101","0101","0100","0100","0110","0101","1000","0011","0001","0001","0001","0001","0101","0111","0100","0011","0011","0101","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1011","0110","0011","0100","0100","0100","0100","0100","0011","0011","0010","0010","0001","0001","0001","0001","0010","0011","0100","0100","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0100","0100","0011","0010","0001","0010","0010","0001","0001","0010","0011","0011","0011","0011","0100","0100","0100","0010","0011","0100","0100","0100","0110","0110","0111","0110","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0100","0110","0110","0100","0100","0011","0100","0100","0101","0101","0101","0110","1011","0111","0111","1000","0011","0011","0010","0010","0011","0011","0010","0011","0011","0011","0011","0010","0011","0100","0110","0110","0110","0110","0110","0111","0111","0110","0101","0100","0101","1001","0101","0000","0010","0110","1011","1100","1011","1011","1011","1011","1011","1010","1011","1011","1010","1011","1100","1011","1011","1100","1100","1010","1011","1011","1011","1000","0101","0101","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0110","0110","0101","0101","0101","1011","1100","1100","0101","1001","1100","1100","1100","1000","0100","0101","0101","0101","0101","0101","0101","0101","0100","1001","1100","1100","1100","1001","0100","0100","1000","1000","0011","0011","0001","0010","0011","0010","0010","0010","0010","0011","0010","0001","0001","0001","0001","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0001","0010","0010","0010","0010","0001","0001","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0010","0010","0010","0010","0001","0001","0010","0010","0010","0001","0010","0011","0010","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1000","1001","1001","1000","1000","0111","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0100","0010","0101","1001","1000","1000","1000","1001","1001","0101","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0100","0100","0011","0011","0011","0100","0100","0100","0011","0010","0001","0001","0010","0011","0100","0010","0010","0100","0011","0100","0101","0100","0100","0100","0101","0101","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0101","0111","0111","1000","1000","1000","1001","1001","1001","1010","1010","1010","0110","0011","0011","0100","0110","1000","1001","1000","1001","1000","1000","1000","1000","1001","1010","1010","1001","1010","1010","1010","1010","1001","1001","1000","1000","1001","1001","1001","1010","1010","1010","1010","1010","1001","0110","0110","0101","0100","0111","0110","1000","0011","0001","0001","0001","0000","0101","0110","0100","0011","0011","0101","1010","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","0101","0011","0011","0100","0011","0011","0011","0100","0100","0011","0010","0001","0001","0001","0001","0010","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0010","0001","0010","0010","0001","0001","0010","0011","0100","0101","0100","0100","0101","0011","0011","0100","0100","0011","0100","0100","0101","0101","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0011","0011","0011","0010","0010","0010","0011","0100","0101","0101","0011","0011","0010","0010","0010","0011","0100","0100","0100","0110","0101","0100","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0110","0100","0100","0110","0111","0110","0111","0110","0110","0110","0110","1000","1010","1011","0101","0010","0100","0111","1011","1010","1010","1011","1010","1010","1010","1010","1011","1010","1011","1011","1011","1011","1100","1011","1000","0111","1010","1011","1011","1010","0100","0011","0011","0011","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0010","0010","0001","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","1011","1100","1100","0110","1001","1100","1100","1100","1000","0100","0101","0101","0101","0101","0101","0100","0100","0100","1001","1100","1100","1100","1001","0100","0011","0011","0100","0100","0011","0100","0100","0100","0011","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0010","0001","0010","0010","0010","0001","0010","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0011","0010","0011","0100","0100","0011","0011","0011","0011","0010","0010","0010","0001","0010","0001","0010","0010","0010","0100","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0100","0100","0111","1000","0101","0110","0100","0010","0011","0011","0010","0011","0011","0010","0010","0010","0100","0010","0101","1001","1000","1000","1000","1000","1000","0100","0010","0010","0011","0010","0100","0011","0010","0010","0010","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","1001","1001","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0010","0010","0010","0011","0011","0011","0011","0100","0100","0010","0010","0100","0101","0011","0001","0010","0100","0100","0100","0100","0011","0000","0001","0011","0011","0100","0010","0010","0100","0010","0011","0100","0101","0100","0100","0011","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0100","0011","0011","0010","0011","0011","0011","0011","0001","0010","0010","0011","0011","0011","0010","0101","0111","0111","1000","1000","1000","1000","1001","1001","1010","1010","1000","0111","0110","0111","0111","0111","1000","1000","1000","1000","1001","1001","1000","1000","1001","1001","1001","1000","1001","1010","1001","1010","1010","1001","1001","1000","1000","1001","1001","1001","1010","1010","1001","1010","1010","1000","0110","0110","0101","1000","0111","1000","0011","0001","0001","0001","0000","0101","0111","0100","0011","0010","0101","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1011","1010","0101","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0001","0010","0100","0100","0100","0100","0100","0011","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0100","0011","0011","0011","0011","0100","0100","0100","0100","0011","0010","0010","0010","0010","0001","0001","0010","0011","0100","0100","0100","0100","0100","0010","0011","0011","0010","0011","0110","0110","0110","0110","0110","0101","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0101","0110","0011","0011","0011","0010","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0001","0100","0100","0011","0100","0101","0101","0101","0101","0101","1000","1001","1010","1010","1001","1000","0111","1000","1001","1010","1010","1010","1010","1010","1011","1011","1010","1010","1011","1011","1011","1011","1100","1011","0101","0001","0001","0011","1010","1100","1011","0101","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0100","0111","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0110","0101","0110","0111","0110","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1011","1100","1100","0110","1001","1100","1100","1100","1001","0101","0101","0101","0101","0101","0100","0100","0100","0100","1001","1100","1100","1100","1001","0100","0100","0100","0100","0100","0100","0100","0101","0101","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0010","0010","0011","0011","0010","0011","0011","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0001","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0100","0100","0100","0100","0011","0011","0010","0010","0001","0010","0010","0001","0001","0001","0010","0101","0110","0110","0110","0110","0110","0101","1000","1000","0100","0101","0110","0111","0110","0111","0110","0101","0101","0100","0011","0011","0010","0011","0011","0010","0010","0010","0101","0011","0101","1001","0111","0111","1000","1000","0111","0100","0010","0010","0011","0010","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","1001","1001","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000"),
("0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0011","0100","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0100","0100","0011","0001","0010","0100","0100","0100","0100","0011","0001","0001","0011","0100","0100","0011","0001","0100","0011","0100","0100","0011","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0010","0011","0011","0010","0010","0001","0001","0010","0011","0011","0011","0010","0101","0111","0111","1000","1000","1000","1001","1001","1001","1001","1001","1000","0111","0111","1000","1000","1000","0111","1000","1000","1000","1001","1001","1001","1001","1000","1001","1000","0111","0100","0100","0100","0100","0100","0100","1000","1001","1001","1000","1001","1001","1001","1001","1000","0101","0100","0101","0110","0111","0011","0100","0101","1000","0011","0001","0001","0000","0000","0100","0111","0100","0011","0011","0101","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","0101","0011","0011","0011","0011","0011","0011","0100","0011","0011","0010","0001","0001","0001","0001","0010","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0010","0001","0010","0010","0001","0001","0001","0001","0011","0100","0011","0101","0011","0010","0011","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0100","0110","0111","0111","0110","0001","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0010","0001","0001","0010","0010","0010","0001","0001","0001","0001","0011","1000","1000","0111","0111","1000","1000","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1000","1001","1010","1000","1001","1010","1001","1001","0100","0000","0001","0101","1010","1000","0110","0101","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0010","0011","0101","0111","0111","0101","0100","0100","0100","0100","0101","0111","1000","1000","1000","0110","0101","1000","1011","1011","1011","1001","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1011","1100","1100","0110","1001","1100","1100","1100","1001","0111","0101","0101","0101","0100","0100","0100","0100","0100","0111","1100","1100","1100","1001","0100","0100","0100","0101","0100","0100","0101","0100","0010","0011","0100","0010","0001","0001","0001","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0011","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0011","0100","0100","0100","0011","0011","0010","0010","0001","0011","0001","0001","0001","0010","0010","0110","0110","0110","0101","0101","0101","0111","1011","0111","0101","0110","1011","1100","1011","1011","1011","1000","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0100","0011","0101","1000","0111","0111","1000","1000","0111","0100","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","1001","1001","1000","0111","1000","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","0111","1000"),
("0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0010","0100","0111","0100","0011","0011","0101","0100","0011","0011","0011","0011","0011","0100","0011","0010","0011","0100","0100","0011","0001","0010","0101","0100","0100","0100","0011","0001","0001","0011","0100","0100","0011","0010","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0001","0001","0001","0010","0010","0011","0011","0011","0101","0111","0111","1000","1000","1000","1000","1001","1001","1001","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1000","1000","1000","0110","0101","0110","0110","0101","0101","1000","1000","1000","1000","1000","1000","1001","1001","1000","0101","0100","0111","1001","1001","0100","0110","0110","0111","0100","0011","0100","0011","0011","0101","0111","0101","0101","0110","0110","0110","0111","0111","1000","0111","0110","0110","0101","1000","1010","1010","1010","1010","1010","0101","0011","0100","0100","0011","0011","0100","0101","0101","0101","0100","0100","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0100","0100","0100","0011","0100","0100","0011","0010","0010","0010","0010","0001","0001","0000","0001","0010","0011","0100","0010","0010","0010","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0011","0100","0100","0101","0110","0101","0110","0110","0110","0110","0110","0101","0110","0110","0101","0101","0111","0111","0111","0101","0100","0100","0101","0110","0011","0011","0010","0010","0011","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","1001","1100","1100","0111","0101","0101","0101","0101","0101","1010","1011","1011","1011","0110","0100","0111","1101","1100","1101","1010","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1011","1100","1100","0110","1001","1100","1100","1100","1000","0100","0100","0101","0101","0101","0100","0100","0100","0100","0011","0111","1011","1100","1001","0011","0011","0011","0100","0011","0011","0100","0011","0010","0011","0100","0010","0010","0010","0010","0010","0001","0001","0001","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0011","0011","0010","0010","0001","0001","0011","0011","0011","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0011","0100","0011","0011","0011","0010","0010","0010","0001","0011","0001","0001","0001","0010","0100","0110","0110","0110","0101","0101","0101","0111","0110","0101","0110","1001","1001","1011","1011","1011","1011","1000","0100","0101","0100","0011","0011","0010","0010","0010","0010","0011","0101","0011","0101","1000","0111","0111","0111","0111","0110","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0100","0110","1001","1001","1000","0111","1000","1000","1000","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","0111","1000"),
("0011","0011","0011","0011","0011","0011","0011","0011","0111","0111","0011","0010","0011","1000","1000","0100","0011","0011","0011","0011","0011","0100","1001","1000","0100","0011","0100","0100","0011","0010","0010","0010","0011","0011","0010","0010","0100","0100","0011","0001","0010","0100","0100","0100","0100","0011","0010","0011","0011","0100","0100","0100","0100","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0100","0011","0001","0001","0000","0001","0001","0010","0011","0011","0011","0101","0111","0111","0111","1000","1000","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1001","1000","0111","1001","0111","0111","0111","0111","0110","0111","1000","0111","1000","1000","1000","1000","1000","1000","0111","0110","0111","1000","0111","0110","1000","0111","1001","1001","1001","1001","1001","1001","1010","1001","1000","1000","1000","1000","1000","0111","0110","1000","1000","1000","1000","1000","1001","1000","1001","1010","1001","1001","1000","0111","0110","0111","1000","1000","1000","1000","1000","1000","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0001","0001","0000","0000","0001","0100","0011","0010","0010","0011","0100","0100","0100","0100","0011","0011","0011","0011","0010","0011","0010","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0100","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0100","0100","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0101","1000","1000","1001","1001","1010","0100","0011","0011","0011","0011","0010","0010","0011","0010","0001","0001","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0011","0100","0100","0100","0101","0101","0101","1010","1100","1100","0111","0101","0101","0101","0101","0101","1010","1010","1011","1100","0110","0100","0111","1100","1100","1100","1010","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1010","1100","1100","0101","1000","1100","1100","1100","1000","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0011","0101","1001","0110","0011","0100","0100","0100","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0010","0001","0010","0010","0010","0011","0011","0011","0011","0011","0100","0101","0101","0011","0001","0010","0010","0010","0011","0101","0110","0110","0100","0010","0010","0010","0100","0101","0100","0011","0011","1001","1011","1011","1011","1000","0100","0100","0100","0100","0100","0011","0010","0010","0011","0101","0101","0011","0110","1000","0110","0111","0101","0110","0110","0100","0101","0101","0100","0100","0011","0010","0010","0100","0101","0101","0101","0101","0101","0100","0100","0101","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0111","1000","1001","1000","0111","1000","1000","1000","1000","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000"),
("0011","0011","0011","0011","0011","0011","0011","0011","0100","1000","1001","0101","0011","0011","0111","1001","0101","0011","0011","0011","0011","0011","0011","0101","0100","0011","0011","0011","0101","0100","0011","0011","0011","0011","0010","0011","0100","0100","0011","0001","0001","0001","0001","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0010","0010","0001","0000","0000","0001","0010","0100","0011","0011","0101","0111","0111","0111","1000","1000","1000","1001","1000","0111","1000","1001","1000","1001","1000","1001","1001","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","0111","0111","1000","1000","0111","1010","1001","0101","0100","0110","0111","0110","0111","0110","0110","1000","1000","1000","0111","1000","0110","1001","1001","0110","0111","0111","0111","1000","0110","0111","1000","1001","1000","1000","1000","1001","1001","1001","1001","0111","1001","1001","0111","1000","1000","0101","0101","0101","0101","0100","0101","0101","0111","1000","0111","0111","0111","1000","1000","1001","1010","1001","1001","1000","1000","1000","1000","1001","0111","0101","0100","0100","0011","0011","0100","0100","0100","0100","0101","0101","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0101","0101","0100","0100","0011","0010","0010","0010","0010","0001","0001","0000","0000","0011","0100","0010","0010","0011","0100","0100","0101","0100","0011","0011","0011","0011","0010","0011","0010","0011","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0101","0011","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0011","0011","0010","0001","0010","0001","0001","0010","0001","0010","0010","0010","0001","0001","0110","1010","1010","1010","1010","1010","0100","0010","0011","0011","0011","0011","0011","0010","0011","0010","0001","0010","0011","0011","0010","0010","0011","0010","0010","0011","1000","1000","0101","0101","0101","0101","0101","0100","1001","1100","1100","0111","0101","0101","0101","0101","0101","1010","1011","1100","1100","0110","0100","0111","1100","1100","1100","1001","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","1010","1100","1100","0110","0011","0111","1100","1100","1000","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0010","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0010","0010","0011","0100","0110","0110","0100","0100","0100","0010","0010","0010","0010","0010","0011","0011","0110","1001","1011","1000","0100","0100","0100","0101","0100","0100","0011","0011","0100","0110","0011","0011","0110","1000","0110","0111","0101","0110","0110","0100","0100","0100","0101","0011","0100","0011","0011","0100","0101","0101","0101","0101","0101","0100","0100","0101","0101","0100","0100","0101","0101","0101","0100","0100","0100","0100","1000","1001","1001","1000","0111","1000","1000","1000","1000","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000"),
("0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0110","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0010","0010","0011","0011","0011","0010","0010","0010","0001","0001","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0010","0001","0000","0000","0000","0001","0011","0011","0011","0011","0101","0111","0111","0111","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","1000","0111","0111","1000","1000","1000","1000","1000","0111","0111","1000","0111","1000","1011","0101","0011","0011","0100","0011","0100","0101","0101","0100","0101","0101","0100","0100","0100","0101","0110","0110","0101","0110","0111","0110","0110","0110","0110","0110","0111","0111","0111","1000","1010","1011","1010","1010","0110","0101","0110","1000","1001","0111","0110","0110","0111","0110","0101","0101","0101","0110","0110","1000","1000","0111","0111","1000","1001","1000","1001","1001","1001","1001","1000","1001","0111","0111","1010","0110","0011","0011","0011","0100","0101","0101","0101","0101","0101","0011","0011","0100","0101","0100","0101","0100","0011","0100","0101","0101","0101","0100","0100","0011","0010","0010","0010","0010","0001","0001","0001","0001","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0011","0100","0010","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0011","0111","0111","0111","0110","0101","1000","1010","1010","1010","1010","1010","0100","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0001","0010","0010","0011","0010","0010","0011","0100","1001","1011","1011","1011","1000","0101","0101","0101","0100","1001","1100","1100","0111","0101","0101","0101","0101","0101","1010","1100","1100","1100","0110","0100","0110","1100","1100","1011","1000","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","1000","1100","1100","0110","0100","0011","0110","1010","0111","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0100","0101","0100","0011","0010","0001","0010","0010","0010","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0010","0010","0010","0001","0011","0011","0010","0010","0011","0011","0011","0100","0101","0011","0001","0010","0011","0010","0100","0110","0010","0011","0110","0100","0101","0110","0110","0100","0011","0011","0011","0011","0100","0100","0011","0100","0111","0111","0100","0100","0100","0100","0100","0011","0011","0011","0100","0110","0100","0010","0110","0111","0100","0100","0011","0011","0010","0100","0100","0101","0101","0011","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0101","1001","1001","1001","1000","0110","1000","1000","1000","1000","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1000"),
("0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0010","0100","0100","0100","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0011","0010","0010","0010","0001","0001","0000","0000","0001","0010","0001","0011","0011","0101","0111","0111","0111","1000","1000","1000","0111","0111","1000","1000","1000","0111","1000","1000","1000","1001","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","1011","0110","0010","0010","0010","0011","0011","0011","0100","0101","0100","0100","0101","0011","0011","0011","0100","0011","0011","0100","0100","0110","0101","0100","0100","0011","0101","0100","0100","0100","0110","0110","0110","0111","1000","0101","0011","0011","0100","0101","0101","0110","1000","1000","0111","0111","0110","0111","0110","0111","1000","1000","1000","1000","1001","0111","0110","0111","1000","1001","1000","1000","0111","0110","1001","1010","1010","0110","0011","0011","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0101","0100","0100","0100","0011","0010","0010","0010","0010","0000","0000","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0011","0010","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0010","0011","0010","0011","0010","0010","0001","0001","0001","0011","1000","1001","0110","1001","1001","1001","1010","1010","1010","1010","1010","1010","0101","0010","0010","0010","0011","0011","0011","0011","0010","0010","0011","0010","0001","0010","0011","0011","0010","0110","1010","1011","1011","1011","1100","1100","1001","0101","0100","0100","1000","1100","1100","0111","0101","0101","0101","0101","0101","1010","1100","1100","1100","0110","0100","0101","0101","1010","1010","1000","1000","0110","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0111","1010","0110","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0010","0001","0010","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0010","0010","0001","0011","0011","0011","0001","0100","0100","0100","0101","1000","0101","0010","0100","0101","0100","0111","1011","0100","0100","0110","0100","0100","0111","0110","0100","0011","0011","0011","0011","0100","0100","0100","0011","0011","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0101","0100","0010","0101","0111","0101","0011","0000","0000","0001","0100","0100","0101","0101","0100","0011","0011","0100","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","1001","1001","1001","1000","0110","0111","1000","1000","1000","1001","1001","1000","1001","1000","1000","1000","1000","1000","1000","1001"),
("0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0011","0011","0011","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0100","0100","0001","0000","0000","0000","0001","0010","0011","0011","0101","0111","0111","0111","0111","1000","1000","0110","1000","1000","1000","0111","0111","1001","0111","1000","1000","0111","1000","1000","1001","1000","1000","1000","1000","1001","0111","1000","0111","0101","1001","1010","0011","0010","0010","0010","0011","0100","0011","0100","0100","0101","0100","0100","0011","0011","0011","0011","0010","0011","0100","0100","0100","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0011","0110","0111","0111","0111","1000","0111","0111","1000","0111","1000","1000","1001","1000","0111","0111","0111","1000","1000","1000","1000","0101","1000","1010","1010","1010","1001","0110","0011","0100","0101","0101","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0001","0010","0010","0010","0010","0011","0100","0100","0100","0100","0101","0011","0100","0011","0011","0011","0010","0010","0010","0100","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0011","0010","0010","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0010","0010","0001","0001","0010","0011","0011","0001","0001","0000","0001","0001","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0010","0010","0001","0011","0111","1000","1001","1000","1000","0111","1000","1001","1010","1010","1010","1010","1010","0101","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0111","1011","1011","1011","1011","1011","1011","1100","0101","0010","0011","0100","0100","1001","1100","0111","0101","0101","0101","0100","0100","0101","1010","1100","1100","0111","0100","0100","0011","0011","1000","1100","1101","1000","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0011","0011","0100","0101","1000","1000","0110","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0010","0010","0001","0010","0011","0011","0010","0011","0100","0100","0101","1001","0110","0011","0101","0100","0100","0110","1010","0100","0100","0101","0101","0100","0110","0110","0100","0011","0100","0011","0011","0011","0100","0100","0100","0011","0100","0100","0100","0101","0101","0101","0101","0101","0100","0101","0101","0100","0011","0101","0111","0101","0011","0001","0000","0001","0100","0100","0101","0101","0100","0100","0011","0011","0100","0100","0100","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0101","1001","1001","1001","0111","0110","0111","1000","1000","1000","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1001"),
("0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0010","0010","0010","0010","0010","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0010","0001","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0001","0000","0000","0000","0000","0010","0011","0011","0010","0100","0111","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","1001","1000","0110","0110","0110","0110","1000","1000","1000","0111","1000","0111","0111","0111","1000","0111","0110","0111","1011","0100","0011","0011","0011","0010","0011","0010","0010","0011","0011","0100","0100","0100","0010","0010","0011","0010","0011","0011","0011","0011","0100","0011","0011","0011","0011","0100","0011","0011","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0100","0110","0111","0111","0111","1000","1000","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","0101","0111","1010","1010","1010","1010","1010","1001","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0011","0010","0011","0011","0010","0010","0010","0011","0100","0010","0010","0010","0001","0001","0001","0001","0001","0010","0010","0011","0010","0010","0011","0011","0010","0100","0101","0100","0011","0011","0011","0011","0010","0001","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0001","0000","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0011","0011","0010","0010","0010","0011","1000","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","0101","0001","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0100","1001","1011","1011","1011","1011","1011","1100","0101","0100","0101","0110","0100","0010","0100","0101","0100","0101","0101","0101","0100","0100","0100","0110","1001","0110","0100","0101","0100","0100","0110","1010","1011","1000","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0110","1100","1101","0111","0100","0101","0101","0101","0101","0100","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0010","0010","0001","0010","0011","0011","0100","0100","0101","0100","0100","0101","0101","0101","0101","0110","0110","0110","0110","0110","0101","0100","0100","0101","0110","0110","0110","0100","0100","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0110","0100","0011","0110","0111","0101","0011","0001","0001","0001","0100","0101","0110","0101","0100","0100","0011","0011","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","1001","1001","1001","0111","0110","0111","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1001"),
("0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0011","0011","0011","0011","0011","0010","0101","1000","0110","0011","0011","0011","0011","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0000","0000","0010","0011","0010","0001","0010","0001","0011","0110","0111","1000","0111","0111","1000","0111","1000","0111","1000","0111","0110","0111","0111","0110","0111","0111","0111","0100","0111","0111","0111","0110","1000","1000","0110","0110","1010","0111","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0100","0011","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0110","0111","1000","1000","1000","1001","1000","1001","1001","1000","1000","1000","1000","1000","1001","0101","0110","1010","1010","1010","1010","1010","1010","1010","1001","0110","0100","0100","0100","0100","0101","0101","0100","0011","0100","0100","0100","0011","0011","0100","0101","0100","0100","0100","0100","0011","0010","0011","0100","0010","0010","0010","0011","0011","0011","0100","0100","0100","0011","0011","0011","0010","0011","0011","0011","0011","0011","0100","0100","0010","0010","0011","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0010","0011","0100","0100","0100","0011","0011","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","0100","0011","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0010","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0001","0100","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0101","0001","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0011","0010","0010","0011","0111","1011","1011","1011","1010","0111","0101","0111","0110","0101","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","1001","1001","0110","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0001","0001","0010","0011","0011","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0010","0010","0010","0010","0001","0001","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0011","0011","0011","0011","0011","0100","0100","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0100","0101","0101","0101","0101","0011","0100","0101","0101","0101","0100","0100","0101","0100","0100","0101","0100","0101","0101","0101","0110","0110","0111","0101","0110","0111","0101","0011","0001","0000","0001","0101","0101","0110","0110","0100","0100","0101","0101","0100","0111","0110","0101","0101","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","1001","1001","1001","0111","0011","0100","0101","0101","0110","1000","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000"),
("0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0111","0100","0010","0011","1000","1000","0100","0011","0011","0011","0011","0011","0101","1001","0101","0010","0010","0011","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0010","0010","0010","0011","0001","0001","0010","0011","0011","0011","0100","0011","0011","0011","0011","0100","0100","0011","0011","0010","0001","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0000","0000","0001","0001","0001","0010","0101","0111","0111","1000","0111","1000","1000","1000","0111","0101","0111","0111","0110","0111","0110","0101","0100","0110","0111","0111","0111","0111","1000","0111","0111","1000","1011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0011","0011","0010","0010","0010","0010","0101","1000","0111","0101","0110","1000","1000","1000","1001","1000","1000","0111","1000","0110","0101","1010","1010","1010","1010","1010","1001","1001","1010","1010","1001","0110","0100","0100","0101","0101","0100","0100","0100","0100","0101","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0011","0011","0100","0100","0011","0011","0010","0010","0010","0010","0011","0010","0011","0100","0100","0100","0011","0010","0010","0010","0010","0001","0000","0000","0001","0001","0001","0010","0010","0010","0011","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0100","0011","0011","0011","0011","0011","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0011","0010","0001","0101","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0101","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0010","0011","0011","0011","0101","1010","0111","0011","0110","0110","0110","0110","0101","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0001","0000","0001","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0001","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0001","0010","0001","0010","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0010","0001","0010","0010","0101","0110","0101","0101","0110","0110","0110","0101","0110","0110","0110","0101","0110","0111","0110","0100","0011","0001","0001","0001","0101","0101","0110","0110","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0101","0011","0011","0100","0101","0101","0111","1000","0101","0010","0010","0011","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0111","1000"),
("0010","0010","0011","0010","0010","0010","0011","0101","0011","0011","0010","0100","1001","0111","0011","0011","0011","0011","0100","1001","1001","0101","0011","0011","1000","1001","0101","0010","0011","0011","0011","0010","0011","0011","0010","0010","0010","0011","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0001","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0010","0010","0011","0010","0010","0011","0011","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0100","0100","0011","0100","0011","0011","0100","0100","0101","0100","0100","0011","0010","0001","0001","0000","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0001","0100","1001","1000","0111","1000","0111","0110","0101","0110","0111","0110","0111","0110","0110","0100","0110","0110","1000","0111","0110","0111","0110","0110","0111","1011","0110","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0100","0100","0011","0011","0100","0011","0100","0011","0011","0101","0100","0011","0010","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0010","0100","0100","0010","0101","1000","0111","0111","0111","1000","0111","1000","0111","0101","1001","1010","1010","1010","1001","1010","1001","1001","1010","1001","1010","1001","0101","0011","0100","0100","0100","0011","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0100","0011","0011","0011","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0000","0000","0000","0000","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0110","1000","0110","0100","0011","0011","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0101","1001","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0110","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0011","0101","0111","0100","0101","0101","0100","0101","0101","0101","0100","0011","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0101","0100","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0010","0001","0010","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0100","0110","0110","0111","0111","0111","0110","0110","0110","0110","0101","0101","0100","0101","0011","0011","0100","0100","0100","0100","0101","0110","0101","0101","0101","0101","0110","1000","0111","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0100","0101","0100","0100","0100","0101","0100","0011","0100","0100","0011","0011","0011","0011","0011","0001","0001","0011","0010","0010","0010","0010","0010","0010","0010","0100","0101"),
("0001","0000","0000","0000","0010","0011","0011","0011","0001","0001","0010","0010","0101","1001","1001","0100","0011","0011","0011","0011","0110","0111","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0001","0001","0010","0011","0011","0101","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0100","0110","0110","0111","0111","0111","0100","0011","0011","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0011","0010","0001","0010","0010","0001","0001","0010","0011","0010","0011","0011","0011","0010","0001","0010","0010","0010","0010","0110","0110","0110","0111","0111","0111","0101","0110","0110","0110","0100","0011","0100","0011","0101","0110","0110","0111","0111","0111","0110","0110","0101","1001","1001","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0001","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0100","1000","1000","0111","1000","1000","1000","1000","0111","0101","1000","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","0101","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0011","0100","0100","0011","0010","0010","0100","0100","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0011","0011","0011","0010","0011","0011","0011","0011","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0110","1001","1001","1001","1010","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0110","0011","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0111","1000","0100","0011","0010","0011","0101","0101","0101","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0100","0010","0010","0010","0100","0100","0100","0101","0101","0101","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0011","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010","0010","0011","0010","0010","0010","0001","0001","0010","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0000","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0011","0010","0010","0010","0001","0010","0100","0100","0011","0011","0100","0011","0011","0100","0011","0100","0101","0110","0100","0011","0100","0100","0100","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0110","0011","0010","0010","0010","0011","0011","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011"),
("0001","0001","0000","0000","0011","0100","0011","0010","0001","0001","0100","0010","0010","0011","0101","0100","0011","0011","0011","0011","0010","0100","0110","0110","0110","0011","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0011","0100","0100","0010","0001","0001","0001","0001","0101","0100","0001","0001","0001","0010","0010","0010","0011","0011","0011","0100","0100","0100","0001","0000","0000","0000","0000","0001","0001","0001","0001","0110","1001","1001","1001","1001","1001","1000","0101","0011","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0011","0101","0100","0100","0011","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0001","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0001","0001","0001","0001","0100","0110","0100","0100","0100","0111","0100","0010","0010","0010","0010","0100","0111","0101","0101","0110","0110","0110","0110","0111","0111","0111","0100","0011","0010","0011","0101","0110","0111","0111","1000","0111","0111","0110","0111","1011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0010","0010","0001","0010","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0100","0110","1000","1000","1000","0111","0111","0100","0110","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1010","1001","0101","0011","0011","0100","0011","0011","0100","0011","0011","0011","0100","0100","0100","0100","0011","0010","0010","0010","0100","0100","0100","0011","0011","0100","0100","0010","0010","0001","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0000","0000","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0001","0001","0001","0010","0010","0011","0011","0010","0001","0001","0010","0010","0010","0001","0001","0010","0010","0001","0010","0010","0010","0011","0111","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0110","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0110","0111","0011","0001","0010","0101","0101","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0001","0010","0010","0011","0101","0101","0100","0101","0100","0100","0010","0010","0011","0011","0001","0010","0011","0011","0011","0010","0001","0001","0001","0001","0000","0001","0001","0001","0001","0010","0001","0001","0001","0001","0011","0010","0001","0001","0010","0010","0100","0100","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0111","0110","0101","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0011","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0001","0010","0001","0001","0001","0001","0001","0010","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0110","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011"),
("0001","0000","0001","0001","0010","0010","0001","0001","0001","0001","0010","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0101","0111","1001","1001","0100","0010","0011","0100","0101","0101","0101","0101","0101","0010","0000","0001","0001","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0101","0101","0100","0101","0110","0111","0111","1000","1000","1000","0111","1000","0111","0110","0010","0001","0001","0001","0001","0001","0001","0001","0010","0101","0111","0110","0110","0110","0101","0101","0101","0011","0011","0011","0011","0100","0100","0100","0011","0011","0001","0010","0011","0011","0101","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0100","0101","0011","0100","0100","0101","0011","0010","0010","0010","0100","0110","0101","0110","0110","0110","0110","0111","0111","0110","0111","0101","0100","0101","0101","0011","0100","0110","0110","0111","0110","0110","0111","0110","1011","0111","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0100","0011","0010","0011","0011","0011","0010","0001","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0010","0101","0111","0111","0111","0101","0101","1001","1001","1001","1001","1001","1010","1001","1001","1001","1001","1001","1001","0111","0110","1001","1010","1001","0101","0011","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0011","0010","0010","0010","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0000","0000","0000","0001","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0100","0100","0010","0010","0010","0011","0011","0011","0011","0010","0001","0001","0010","0010","0001","0010","0001","0010","0010","0010","0001","0010","0011","1000","1010","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","1010","1010","1010","1000","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0100","0100","0010","0010","0011","0101","0101","0100","0100","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0101","0101","0100","0101","0101","0101","0100","0100","0100","0100","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0010","0010","0011","0011","0101","0101","0101","0101","0100","0100","0100","0100","0101","0100","0011","0010","0011","0100","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0101","0100","0011","0111","1001","1000","1000","1000","1000","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1001","1010","1001","1000","1000","1000","0110","0110","0100","0101","0011","0101","0100","0101","0110","0100","0011","0010","0011","0011","0011","0100","0101","0011","0101","0101","0100","0100","0011","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0101","0101","0001","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0001","0000","0000","0001","0000","0001","0001","0001","0001","0001","0001","0001","0100","0111","0111","0110","0010","0010","0011","0011","0011","0110","0111","0110","1000","0100","0010","0100","0101","0101","0110","0110","0110","0110","0011","0000","0001","0001","0010","0011","0001","0000","0010","0011","0001","0001","0001","0001","0100","1000","1000","0111","1000","0111","0111","0111","0111","0110","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0100","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0011","0011","0010","0010","0010","0011","0101","0101","0101","0110","0110","0101","0101","0110","0110","0111","0110","0101","0101","0110","0101","0011","0100","0110","0110","0110","0110","0110","0110","1000","1010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0011","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0111","1000","0101","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0100","0011","1000","1001","1010","1001","0101","0100","0100","0011","0100","0011","0100","0100","0100","0100","0011","0011","0010","0010","0011","0101","0100","0100","0100","0101","0100","0011","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0000","0000","0000","0000","0001","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0011","0010","0010","0010","0010","0011","0011","0011","0010","0001","0001","0001","0001","0001","0010","0001","0010","0011","0010","0010","0011","1000","1010","1001","1010","1010","1010","1001","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1011","1010","1010","1010","1000","0011","0011","0011","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0100","0101","0101","0100","0011","0010","0011","0100","0100","0001","0001","0001","0001","0001","0001","0010","0100","0100","0100","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0010","0001","0010","0010","0100","0100","0010","0010","0111","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","1000","1000","1001","1000","0110","0111","0110","0101","0100","0101","0101","0100","0011","0100","0011","0011","0100","0010","0010","0010","0100","0100","0011","0100","0100","0011","0101","0110","0101","0101","1000","0110","0100","0101","0101","0011","0010","0010","0001","0001","0001","0010","0010","0010","0010","0001","0001","0001","0000","0001","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0010","0010","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0110","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0011","0100","0100","0110","0111","0111","0010","0010","0100","0101","0101","0110","0111","0111","0110","0111","0111","0101","0101","1000","1000","1000","0111","0111","0011","0001","0001","0001","0101","0110","0010","0001","0011","0011","0010","0010","0010","0010","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0011","0100","0011","0010","0010","0010","0010","0011","0100","0100","0101","0101","0100","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0011","0100","0100","0011","0010","0011","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0010","0011","0011","0100","0111","1010","1011","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0110","0011","1001","1001","1001","1001","1001","0110","0011","0011","0100","0100","0100","0100","0011","0010","0010","0010","0011","0011","0011","0010","0010","0010","0100","0100","0100","0011","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0000","0001","0001","0000","0000","0000","0000","0000","0001","0001","0010","0010","0011","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0001","0001","0001","0010","0010","0010","0010","0010","0000","0001","0001","0001","0010","0001","0001","0010","0010","0010","0100","1000","1010","1001","1010","1010","1010","1010","1001","1001","1010","1011","1011","1010","1010","1011","1011","1010","1010","1011","1011","1011","1011","1010","1010","1010","0111","0010","0100","0100","0011","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0001","0010","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0001","0001","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0011","0011","0011","0010","0001","0001","0001","0100","0100","0001","0001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1001","1001","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0101","0101","0101","0101","0101","0101","0100","0011","0010","0010","0010","0011","0100","0011","0011","0011","0100","0011","0010","0100","0100","0011","0011","0101","0101","0101","0110","0110","0100","0110","0111","0110","0110","0101","0101","0110","0111","0110","0101","0101","0100","0011","0010","0001","0001","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0001","0010","0010","0001","0010","0010","0010","0010","0001","0010","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010"),
("0010","0010","0000","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0111","0111","0111","1000","1000","0111","0110","1001","1001","1000","1000","0111","0100","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0010","0011","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0011","0100","0011","0010","0010","0011","0100","0011","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0001","0011","0010","0011","0010","0010","0010","0011","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010","0011","0011","0011","0010","0010","0101","0110","0110","0111","1001","1001","1001","1001","1001","1000","1001","1001","1000","1001","0110","0100","1000","1001","1001","1001","0111","0101","0011","0100","0100","0100","0100","0011","0010","0010","0011","0011","0100","0011","0010","0010","0011","0100","0100","0100","0100","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0001","0000","0000","0001","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0001","0001","0001","0001","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0001","0010","0010","0010","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1010","1010","1011","1011","1010","1010","1010","1010","1011","1010","1010","1010","1010","1010","0110","0010","0011","0011","0010","0001","0001","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0010","0010","0011","0110","0101","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0011","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","0111","0110","0111","0111","0111","1001","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0110","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0101","0100","0101","0100","0100","0011","0010","0011","0011","0010","0011","0100","0100","0101","0100","0010","0010","0011","0110","0011","0010","0010","0100","0100","0101","0110","0110","0100","0101","0110","0101","0101","0101","0111","0111","0111","0111","0110","0100","0110","0011","0010","0010","0011","0010","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0001","0001","0001","0010","0010","0010","0010","0001","0010","0001","0010","0010","0010","0001","0001","0010","0010","0001","0010","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0101","0101","0010","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0010","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0000","0001","0010","0001","0001","0000","0011","0111","0110","0111","1000","1000","1000","0110","1001","1000","0111","0101","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0001","0010","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0011","0010","0010","0010","0010","0100","0010","0010","0011","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0010","0011","0010","0011","0011","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0010","0010","0011","0011","0101","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0110","0100","1001","1001","0111","0100","0011","0100","0100","0100","0100","0100","0010","0010","0010","0011","0100","0100","0011","0010","0011","0100","0100","0100","0100","0100","0010","0001","0001","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0001","0001","0000","0000","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0100","0100","0011","0011","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0010","0101","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0110","0010","0100","0100","0010","0010","0010","0100","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0100","0101","0100","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0111","0011","0010","0010","0010","0010","0100","0111","1000","1001","1000","1000","1000","0111","0110","0110","0101","0101","0100","0100","0100","0100","0110","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0101","0110","0101","0111","1000","1000","1000","0111","1000","0110","0110","0111","0110","0110","0111","0110","0100","0101","0110","0101","0011","0011","0011","0010","0010","0010","0010","0011","0100","0011","0011","0011","0010","0100","0011","0011","0010","0011","0011","0011","0100","0100","0011","0100","0100","0011","0011","0101","0110","0101","0100","0101","0101","0101","0110","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0110","0100","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010"),
("0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0001","0001","0000","0001","0010","0001","0001","0001","0010","0111","1000","0111","1000","1000","1000","0110","1000","0101","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0100","0011","0011","0011","0001","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0011","0011","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0011","0010","0011","0011","0100","0100","0101","1000","1001","1001","1001","1001","1001","1000","1001","1000","1001","0111","0100","0111","0101","0100","0100","0100","0100","0100","0100","0100","0010","0001","0010","0010","0011","0011","0011","0100","0011","0011","0011","0100","0100","0100","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0010","0010","0001","0001","0001","0000","0000","0000","0001","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0101","0110","0111","0111","0110","0101","0101","0101","0101","0110","0111","0110","0111","0111","0111","0111","0110","0111","0110","0110","0110","1000","1000","0111","0111","0111","1000","1000","1001","1001","1001","1001","1001","1010","1001","1010","1001","1010","1010","1011","1010","1010","1010","1010","1011","1011","1010","1010","1011","1011","1011","1011","0110","0010","0011","0011","0010","0001","0001","0010","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0100","0001","0010","0010","0010","0101","0101","1000","1000","1001","1001","0110","0001","0001","0001","0010","0010","0010","0001","0001","0001","0101","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0101","0101","0100","0101","1000","1000","0111","0110","0111","0110","0111","0110","0101","0100","0100","0110","0110","0100","0100","0101","0100","0010","0011","0011","0010","0100","0010","0010","0010","0010","0100","0100","0011","0010","0100","0011","0010","0100","0010","0011","0011","0100","0011","0011","0010","0010","0100","0101","0110","0110","0100","0100","0101","0101","0110","0011","0011","0010","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0001","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0001","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0010","0010","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0011","0111","0011","0011","0011","0010","0010","0011","0011","0011","0010","0011","0010","0010","0010","0001","0010","0001","0001","0010","0010","0010","0011","0010","0010"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0110","0110","0111","0111","0111","0101","0011","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0011","0011","0011","0010","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0010","0011","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0100","0100","0011","0011","0110","1001","1001","1000","1000","1000","1000","1000","1000","0110","0011","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0011","0010","0010","0010","0100","0100","0100","0100","0100","0100","0100","0011","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0000","0001","0011","0011","0011","0011","0100","0100","0001","0001","0010","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0100","0100","0110","0111","1000","1000","1000","0111","0111","0110","0110","0110","0101","0110","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","1000","0111","0111","0111","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1001","0101","0011","0100","0100","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0001","0011","0010","0001","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0101","0011","0011","0011","0011","0110","0110","1000","1000","1001","1001","0111","0010","0010","0010","0001","0001","0001","0010","0001","0010","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0110","0111","0110","0100","0011","0100","0101","0101","0101","0101","0101","0110","0110","0110","0110","0100","0100","0100","0100","0010","0011","0100","0011","0010","0011","0011","0010","0011","0011","0011","0010","0010","0011","0100","0011","0010","0011","0011","0010","0010","0010","0100","0100","0100","0100","0011","0011","0011","0110","0101","0101","0100","0011","0101","0111","0110","0111","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0001","0001","0010","0011","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0100","0101","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0001","0001","0000","0001","0010","0010","0011","0010","0010"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0011","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0100","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0001","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0001","0010","0010","0010","0001","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0011","0100","0100","0011","0010","0010","0100","1000","1001","1000","1000","1000","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0011","0011","0010","0010","0010","0011","0100","0100","0100","0100","0101","0100","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0000","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0101","0110","0111","0101","0001","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0101","0111","0111","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0111","0111","0111","0110","0110","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0110","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0111","0111","0111","1000","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0101","0011","0011","0010","0011","0110","0110","1000","1001","1001","1000","1000","0011","0011","0011","0010","0010","0010","0010","0010","0010","0110","1000","0111","1000","1000","1001","1001","1000","1000","1000","1000","1000","0111","0101","0101","0110","0101","0100","0010","0011","0101","0011","0100","0110","0100","0100","0101","0101","0100","0100","0110","0101","0011","0100","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0010","0100","0011","0001","0010","0010","0010","0011","0101","0101","0100","0101","0100","0011","0101","0100","0100","0011","0100","0101","0101","0111","0111","0100","0011","0011","0011","0010","0011","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0001","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0001","0010"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0100","0100","0011","0011","0010","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0011","0011","0011","0011","0100","0100","0011","0011","0100","0011","0100","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0010","0010","0010","0001","0001","0010","0010","0001","0001","0100","0011","0011","0100","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0100","0100","0011","0010","0010","0010","0100","0110","1000","0110","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0010","0100","0100","0100","0100","0100","0100","0011","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0000","0000","0000","0001","0010","0011","0010","0011","0011","0011","0111","1001","1011","1100","1101","1101","1101","1100","1001","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","1000","0111","0111","1000","0111","1000","0111","0111","1000","0111","1000","0111","0111","1000","1000","1001","1000","1000","1000","1000","1001","1000","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0110","0110","0110","0101","0101","0101","0101","0100","0100","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0011","0010","0011","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0101","0010","0011","0010","0011","0110","0110","1000","1001","1001","1001","1000","0100","0011","0011","0011","0010","0010","0010","0010","0001","0110","1000","0111","0111","1000","1001","1000","1000","1000","1000","1000","1000","1000","0111","0111","0110","0110","0100","0100","0011","0011","0011","0101","0110","0101","0100","0100","0100","0011","0011","0011","0100","0011","0011","0010","0001","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0010","0001","0001","0001","0011","0100","0110","0111","0101","0100","0100","0100","0101","0101","0010","0011","0101","0101","0110","0101","0111","0100","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0011","0010","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0001","0001","0010","0001","0001","0001","0010","0010","0010","0001","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0001","0001","0001","0010","0010","0001","0010"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0011","0011","0100","0100","0011","0011","0010","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0110","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0001","0001","0001","0001","0001","0010","0010","0010","0001","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0010","0010","0100","0101","0010","0010","0010","0001","0010","0010","0010","0001","0010","1010","1000","0111","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0001","0011","0001","0010","0010","0001","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0100","0100","0100","0010","0010","0010","0010","0010","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0100","0100","0010","0010","0010","0010","0001","0010","0100","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","1000","1001","1011","0110","0010","0010","0010","0011","0100","0111","0111","1100","1101","1101","1101","1101","1101","1101","1101","1001","0011","0011","0101","0110","0110","0100","0010","0010","0011","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0110","0111","0111","0110","1000","0110","0111","1000","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","1000","0111","0111","0111","1000","1001","0111","1000","0111","0111","1000","0111","0111","0111","0110","0111","0111","0111","1000","0111","1000","0111","0111","1000","0111","1000","0111","0111","0100","0011","0011","0011","0010","0101","0101","0110","0110","0110","0110","0110","0111","0110","0101","0110","0111","1000","1000","1000","1000","0111","0111","0111","0111","1000","0111","0101","0100","0100","0011","0011","0110","0110","1000","1000","1000","1000","0111","0010","0001","0010","0010","0001","0001","0001","0001","0001","0101","1000","0111","0111","1001","1001","1000","1000","1000","1001","1001","1000","0111","0111","0111","0110","0111","0110","0100","0100","0011","0100","0101","0101","0100","0101","0011","0100","0011","0011","0010","0010","0010","0010","0010","0001","0001","0100","0100","0011","0010","0001","0010","0001","0010","0011","0010","0011","0010","0010","0011","0010","0010","0010","0011","0100","0101","0110","0110","0100","0101","0011","0101","0100","0011","0100","0100","0011","0100","0101","0101","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0001","0010","0010","0010","0001","0001","0010","0001","0001","0001","0001","0010","0001","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0101","0011","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0010","0001","0001","0001","0010","0010","0001","0001","0010","0010","0010","0001","0001","0010","0001","0100","0100","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001"),
("0010","0010","0010","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0011","0011","0010","0010","0011","0100","0100","0100","0011","0100","0100","0010","0010","0010","0001","0010","0010","0001","0001","0011","0110","0111","0101","0010","0001","0010","0010","0100","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0100","0100","0100","0010","0001","0010","0001","0001","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0111","1010","1011","1011","0110","0010","0010","0010","0011","0100","1000","1001","1101","1101","1101","1101","1100","1011","1010","1001","1000","0111","0111","0111","0111","0110","0110","0100","0010","0011","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0110","0110","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","1000","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0111","1000","1000","0111","1000","0111","1000","0111","0111","1000","0110","0111","0111","0111","1000","0111","0111","0111","0111","1000","0111","0111","1000","0111","0110","0011","0011","0011","0011","0101","0110","0110","0110","0110","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","0111","1000","0111","0111","0111","0110","0111","0111","1000","1000","0111","0110","0111","0111","0111","0110","0110","0110","0110","0110","0010","0000","0001","0001","0010","0010","0010","0001","0001","0101","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0110","0110","0110","0100","0100","0100","0011","0100","0100","0100","0100","0010","0010","0010","0011","0011","0010","0011","0010","0011","0010","0001","0011","0011","0010","0010","0010","0001","0001","0011","0011","0011","0010","0010","0010","0011","0011","0001","0010","0011","0100","0100","0101","0101","0100","0110","0101","0100","0011","0011","0110","0110","0110","0101","0110","0110","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0010","0010","0001","0010","0011","0100","0010","0010","0010","0010","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0011","0001","0001","0001","0011","0011","0011","0010","0100","0101","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0001","0001","0010","0010","0010","0010","0010","0010","0011","0010","0001","0010","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0011","0010","0010","0011","0011","0011","0010","0101","1010","1001","0111","0110","0110","0110","0110","0101","0100","0011","0100","1000","1011","1001","0110","0101","0101","0101","0101","0100","0011","0010","0010","0010","0010","0001","0001","0001","0010","0001","0001","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0111","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0010","0001","0001","0010","0010","0001","0001","0010","0010","0010","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0100","1000","1001","1100","1011","1010","1001","0111","0111","0110","0110","0110","0110","0111","0111","0111","0111","0110","0110","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0111","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0111","0111","0110","0111","1000","0110","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","1000","0110","0111","0111","0110","0111","0111","1000","1000","0111","0111","0111","0111","0111","0110","0111","0111","0111","1000","0111","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","0111","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0111","0111","0111","1000","1000","1000","1000","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0111","1000","0110","0111","0110","0110","0111","0011","0001","0010","0010","0010","0010","0010","0010","0010","0101","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","1000","0111","0101","0101","0101","0011","0010","0010","0011","0100","0011","0011","0010","0010","0010","0010","0011","0010","0011","0011","0011","0011","0010","0010","0010","0001","0001","0010","0001","0010","0011","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0110","0110","0011","0010","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0001","0010","0001","0001","0010","0001","0010","0010","0001","0001","0000","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0010","0010","0010","0011","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0000","0000","0001","0001","0001","0011","0011","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0100","0001","0001","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0110","1000","1000","0101","0100","0100","0110","0111","0101","0100","0110","0110","0110","0110","0110","0101","0100","0100","0101","0101","0100","0101","0110","0110","0110","0110","0101","0100","0100","0011","0011","0010","0001","0010","0010","0001","0001","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","1000","0100","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0010","0001","0001","0010","0010","0001","0001","0010","0010","0010","0011","0100","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0100","0111","0111","0111","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0110","0111","1000","0111","0111","0110","0111","0110","0110","0110","0110","0111","0110","0110","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","1000","0111","0111","0111","0111","1000","0110","0111","0111","0110","0111","0111","0111","1000","0111","1000","0111","0111","0111","0110","0111","1000","1000","0111","0110","0111","0111","0110","0111","0111","0110","0110","0110","0110","0110","0110","0111","0111","1000","1000","0111","1000","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","1000","0111","0111","0111","0111","1000","0111","0110","0111","0110","0111","0110","0011","0010","0011","0011","0010","0010","0010","0010","0010","0110","1000","0111","1000","1000","1000","1000","1000","0111","1000","0111","0111","0111","1000","1000","0111","0101","0100","0011","0011","0010","0010","0011","0011","0011","0011","0010","0011","0100","0101","0101","0100","0011","0011","0010","0010","0001","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0011","0011","0011","0010","0101","0101","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0010","0001","0001","0001","0001","0001","0010","0001"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0011","0010","0001","0000","0000","0000","0001","0000","0001","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0010","0011","0011","0010","0010","0010","0001","0001","0001","0000","0001","0001","0001","0011","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0100","0011","0100","0011","0011","0011","0100","0100","0101","0101","0100","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0001","0010","0011","0111","1000","0110","0101","0110","0110","0110","0100","0101","0100","0110","1000","0111","0101","0101","0101","0100","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0011","0100","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0011","0011","0010","0010","0001","0001","0001","0001","0000","0000","0001","0010","0010","0010","0010","0010","0010","0011","0100","0101","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0100","0010","0001","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0101","1010","1011","1100","1101","1010","0011","0001","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0100","0101","0110","0110","0101","0110","0111","0111","0110","0110","0111","0111","0111","0111","0110","0110","0110","0110","0110","0111","0110","0111","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0101","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0111","0110","0110","0111","0110","0111","0110","0110","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","1000","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0111","1000","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","1000","0111","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0111","1000","0110","0110","0110","0110","0110","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0110","0111","0110","1000","0111","0110","0111","0110","0110","0111","0101","0100","0010","0011","0010","0010","0010","0010","0010","0010","0101","1001","1000","1000","1001","1000","1001","1000","0110","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0100","0011","0011","0010","0010","0010","0011","0010","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0011","0011","0010","0010","0010","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0010","0011","0100","0011","0010","0011","0100","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001"),
("0001","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0101","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0011","0001","0001","0001","0001","0001","0001","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0011","0010","0010","0001","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0011","0100","0101","0011","0001","0001","0001","0010","0010","0010","0010","0010","0110","1000","0111","0100","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0101","0101","0101","0100","0101","0100","0101","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0100","0011","0011","0010","0010","0010","0010","0000","0001","0011","0011","1000","0100","0011","0010","0010","0011","0101","0101","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0101","0100","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0010","0011","0011","0011","0101","1000","0111","0100","0101","1001","1100","1000","0010","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0010","0011","0100","0101","0110","0111","0111","0111","0111","0111","0110","0111","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","1000","1000","0111","1000","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","1000","1000","0111","0111","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","1000","0111","0110","0110","0110","0111","0110","0110","0111","0111","1000","0111","0111","1000","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","1000","0110","0111","0110","0111","1000","0111","0111","0111","0110","0111","0110","0110","0011","0010","0011","0011","0010","0010","0010","0010","0010","0100","1000","0111","1000","1001","1001","1001","1000","0110","0010","0010","0001","0010","0010","0010","0010","0001","0011","0011","0011","0010","0010","0011","0010","0011","0100","0011","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0010","0010","0001","0000","0001","0001","0000","0001","0001","0001","0010","0001","0010","0010","0010","0010","0010","0001","0000","0011","0001","0010","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0001","0011","0101","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010"),
("0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0100","0101","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0100","0011","0011","0011","0011","0010","0010","0010","0001","0000","0000","0000","0000","0000","0001","0010","0011","0100","0010","0010","0001","0010","0010","0011","0011","0011","0100","0011","0010","0010","0011","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0100","0110","0110","0101","0101","0101","0100","0100","0011","0010","0010","0010","0011","0011","0011","0100","0110","0011","0100","0100","0100","0100","0011","0011","0100","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0010","0010","0011","0100","0111","1000","0101","0011","0101","0110","0110","1010","1001","0010","0001","0010","0001","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0011","0100","0110","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0110","0011","0100","0110","0111","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","1000","1000","1000","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","1000","0111","0111","0111","0111","1000","0111","0110","0111","0110","0110","0110","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","1000","0111","0111","0111","0111","1000","0111","0110","0111","0110","0111","0111","0110","0110","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0101","0111","1000","1001","1001","1001","1000","0111","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0001","0010","0011","0100","0010","0011","0001","0001","0001","0001","0010","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0010","0011","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0001","0001","0010","0010","0000","0001","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0001","0001","0100","0110","0010","0001","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010"),
("0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0101","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0011","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0101","0110","0101","0101","0100","0011","0010","0100","0011","0111","0011","0011","0100","0110","0101","0100","0100","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0101","0101","0101","0101","0101","0011","0100","0011","0010","0010","0011","0011","0011","0011","0100","0111","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0010","0010","0001","0001","0100","0101","0101","0101","0011","0100","0101","0101","0101","0101","0100","0101","0101","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0101","0101","0100","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0010","0010","0001","0010","0011","0101","1000","0111","0100","0011","0010","0010","0100","0100","0110","0110","0011","0010","0001","0001","0010","0001","0010","0010","0010","0011","0010","0001","0001","0001","0010","0011","0101","0110","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0110","0101","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0111","0100","0100","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0111","1000","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0110","0111","1000","0110","0111","0111","0111","0111","0111","1000","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","1000","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","1000","0111","0110","0111","0110","0111","0111","0110","0111","0111","0110","0111","0110","0111","0110","0110","0110","0101","0101","0100","0011","0011","0100","0100","0100","0011","0101","1000","1001","1001","1001","1000","0111","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0010","0001","0010","0010","0010","0010","0011","0001","0001","0001","0001","0010","0001","0001","0001","0001","0011","0011","0011","0011","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0010","0010","0011","0010","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0101","0111","0100","0010","0010","0001","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010"),
("0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0101","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0101","0101","0101","0101","0101","0100","0011","0011","0101","0111","0011","0010","0101","0110","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0101","0101","0101","0101","0100","0011","0100","0011","0010","0010","0010","0011","0011","0011","0011","0110","0100","0000","0000","0000","0000","0000","0001","0011","0011","0011","0011","0011","0010","0001","0010","0010","0011","0011","0010","0010","0011","0100","0101","0110","0110","0110","0101","0101","0100","0011","0010","0010","0010","0010","0010","0010","0001","0010","0100","0101","0100","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0010","0010","0011","0100","0110","1000","1000","1100","1010","0011","0011","0011","0011","0001","0010","0011","0101","0110","0011","0010","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0101","0110","0111","1000","1000","1000","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0110","0110","0110","0111","0110","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0110","0101","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0100","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","1000","0111","1000","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","1000","0111","0111","0111","0110","0111","0111","0111","1000","0111","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","1000","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","1000","1000","0110","0111","0110","0111","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0100","0011","0111","1001","1001","1001","1000","0110","0011","0100","0100","0011","0010","0010","0001","0001","0001","0010","0010","0010","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","0011","0100","0011","0010","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0010","0010","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0110","0111","0110","0010","0010","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0100","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0100","0011"),
("0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0101","0011","0011","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0100","0100","0100","0100","0100","0011","0100","0001","0010","0010","0010","0010","0010","0010","0001","0001","0001","0000","0000","0000","0000","0000","0001","0011","0011","0011","0011","0011","0011","0011","0001","0000","0001","0010","0101","0100","0101","0101","0101","0110","0110","0110","0110","0110","0101","0100","0100","0011","0011","0011","0010","0010","0001","0010","0100","1001","1010","0011","0001","0001","0001","0010","0100","0100","0100","0100","0100","0100","0111","1000","1001","1000","1000","0111","0101","0110","0101","0011","0011","0011","0010","0010","0010","0011","0011","0100","0010","0001","0001","0001","0010","0010","0010","0010","0011","0011","0100","0111","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0101","0101","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0111","1001","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0111","0111","0101","0011","0101","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0111","1000","0110","0110","0111","0111","0111","0110","0110","0111","0111","1000","0111","0110","0111","0110","1000","1000","0111","0111","0111","0111","1000","0110","0111","0111","0111","1000","0111","0111","1000","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0111","0111","0110","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","1000","1001","1001","0111","0110","0101","0101","0101","0100","0010","0001","0010","0010","0101","0100","0010","0010","0001","0001","0001","0001","0010","0011","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0100","0100","0100","0100","0011","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0100","0111","0111","0110","0011","0010","0010","0010","0010","0001","0010","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0100","0101","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0011","0011","0010","0010","0011","0011","0011","0011","0010","0011","0110","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0011","0010","0010","0001","0001","0001","0001","0010","0001","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0011","0010","0010","0011","0011","0011","0011","0100","0101","0101","0100","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0100","0100","0010","0010","0001","0011","0100","0110","1010","0111","0110","0111","0110","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0100","0101","0101","0100","0101","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0110","0111","0111","0111","0111","0111","0110","0110","0110","0110","0111","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0111","1000","1000","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0110","0110","0111","0110","0110","0111","0110","0111","0111","0111","0111","0110","1000","1000","0111","0111","0111","0101","0100","0110","0111","0111","0110","0111","0111","1000","0111","0110","0111","0111","0111","0111","0110","0110","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","1000","0111","0111","1000","0101","0100","0111","0111","0111","0110","0111","0111","0110","0111","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","1001","0111","0101","0101","0101","0101","0100","0101","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0101","0100","0010","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0011","0010","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0011","0010","0010","0101","0111","0111","0111","0101","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010"),
("0010","0011","0011","0010","0001","0010","0010","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0100","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0101","0101","0011","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","0111","0101","0101","0110","0110","0101","0011","0011","0101","0101","0101","0101","0100","0100","0100","0100","0100","0010","0010","0011","0100","0011","0011","0011","0011","0010","0010","0011","0011","0100","0100","0101","0110","0110","0110","0101","0100","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0011","0010","0011","0100","0011","0100","0110","0111","0110","0100","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0100","0100","0100","0100","0101","0011","0001","0001","0001","0001","0010","0101","0110","0101","0101","0100","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0110","1000","0111","0111","0111","0111","1000","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0101","0011","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0110","0111","0111","0110","0101","0110","0111","0111","0110","0111","0110","0111","0111","0110","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0111","1000","0101","0101","0100","0100","0100","0100","0011","0010","0010","0010","0011","0010","0010","0001","0001","0001","0010","0001","0001","0010","0001","0001","0001","0001","0010","0001","0001","0001","0010","0100","0011","0100","0011","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0011","0010","0011","0010","0010","0010","0011","0100","0100","0100","0100","0011","0011","0011","0011","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0001","0010","0110","0111","0111","0111","0110","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0010"),
("0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0011","0110","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","1000","0110","0010","0100","1000","1000","0110","0010","0011","0110","1000","1000","1000","1000","1000","0111","0111","0111","0011","0010","0100","0110","0101","0011","0011","0010","0011","0011","0011","0011","0011","0100","0101","0101","0110","0110","0110","0110","0101","0011","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0100","0011","0010","0011","0011","0011","0011","0011","0001","0010","0001","0010","0010","0001","0010","0001","0011","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0110","0100","0001","0001","0001","0001","0001","0010","0011","0100","0101","0101","0011","0011","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0111","0111","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","1000","1000","0110","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0110","0111","0111","0111","1000","0111","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0101","0110","0110","0110","0110","0101","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0010","0010","0011","0011","0010","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0010","0010","0010","0011","0011","0011","0010","0010","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0100","0110","0111","0111","0110","0110","0100","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0010"),
("0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0011","0010","0100","0100","0100","0100","0100","0100","0101","0011","0000","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0101","0110","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1000","0111","0011","0100","0111","1000","0110","0010","0010","0110","0111","0111","1000","1000","1000","1000","0111","0111","0101","0101","0101","0101","0101","0101","0100","0010","0010","0010","0010","0011","0011","0100","0101","0101","0101","0110","0110","0110","0110","0101","0100","0011","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0100","0010","0010","0010","0010","0010","0011","0010","0011","0010","0100","0100","0011","0100","0011","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0110","1000","1001","0110","0010","0001","0001","0001","0001","0001","0010","0010","0100","0101","0101","0101","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0111","1000","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0111","1000","0110","0111","0110","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","1000","0111","0111","1000","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0110","0110","0011","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0100","0010","0010","0011","0100","0011","0011","0010","0001","0010","0010","0010","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0010","0011","0010","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0101","0111","0110","0111","0111","0111","0101","0010","0010","0010","0011","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010"),
("0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","0011","0101","0101","0101","0101","0101","0101","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0011","0110","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","1000","0101","0110","0111","0111","0111","0100","0101","0110","0111","0111","0111","0111","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0010","0010","0010","0011","0100","0100","0101","0101","0110","0110","0110","0110","0101","0110","0110","0100","0011","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0100","0100","0100","0100","0100","0011","0100","0010","0100","0011","0011","0100","0011","0101","0101","0100","0100","0101","0101","0110","1000","1000","1001","1010","1001","0111","0010","0001","0001","0001","0001","0001","0001","0001","0010","0011","0101","0110","0111","0111","0110","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","1000","1000","0111","0111","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0110","1000","0110","0110","0111","0111","1000","0111","0110","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0101","0011","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0100","0011","0010","0011","0011","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0100","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0011","0100","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0011","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0110","0111","0110","0111","0111","0111","0110","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0001","0010","0011","0010","0011","0011","0010","0010"),
("0110","0110","0101","0101","0101","0101","0101","0101","0101","0110","0101","0011","0101","0110","0110","0110","0110","0101","0011","0001","0001","0010","0010","0010","0010","0010","0100","0110","0101","0010","0100","0110","0011","0011","0101","0011","0010","0101","0100","0010","0011","0011","0010","0011","0011","0010","0010","0011","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0100","1000","1000","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","1000","0101","0110","1000","1000","0111","0100","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0010","0010","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0011","0011","0101","0110","0110","0110","0110","0101","0110","0110","0110","0101","0101","0101","0101","0101","0100","0100","0100","0011","0100","0010","0100","0101","0011","0100","0011","0100","0101","0110","1000","1010","1010","1011","1011","1011","1010","1010","1000","0011","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0110","0110","0101","0101","0111","0110","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","1000","0111","0111","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0111","0111","1000","0110","0111","0111","0101","0111","0111","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0111","1000","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0110","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0100","0100","0010","0011","0011","0010","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0001","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0100","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0100","0110","0111","0111","0111","0110","0111","0110","0100","0000","0000","0000","0000","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0010","0010","0010","0010","0010","0010"),
("0101","0100","0011","0010","0011","0011","0011","0011","0011","0100","0011","0011","0110","0110","0110","0110","0110","0101","0001","0001","0010","0010","0010","0010","0010","0011","0110","1000","0100","0011","0111","0111","0011","0110","0111","0011","0101","1000","0100","0100","0111","0011","0100","0111","0110","0010","0101","0111","0100","0011","0110","0101","0010","0110","0101","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0010","0100","0011","0010","0011","0011","0010","0011","0011","0011","0010","0011","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0010","0011","0010","0011","0011","0011","0011","0011","0010","0011","0110","0110","0100","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","1001","0110","0110","0111","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0011","0011","0101","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0100","0011","0100","0100","0010","0010","0100","1001","1011","1100","1100","1100","1011","1010","1011","1011","1010","1001","0011","0001","0001","0001","0001","0001","0010","0010","0011","0010","0001","0100","0110","0101","0100","0011","0101","0110","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0110","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0111","1000","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0111","1000","0111","0111","1000","0110","0110","0110","0111","1000","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0110","0111","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0101","0111","0110","0111","0110","0110","0110","0110","0101","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001"),
("0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0110","0111","0111","0110","0110","0011","0001","0010","0010","0010","0010","0010","0010","0101","1000","0110","0010","0110","1000","0100","0100","1000","0101","0011","1000","0111","0011","0110","0101","0011","0111","1000","0101","0011","0111","0111","0011","0110","1000","0100","0101","0110","0011","0011","0011","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0011","0011","0101","1000","0101","0011","0111","0111","0010","0110","0111","0011","0101","0101","0010","0011","0110","0100","0010","0110","0100","0010","0101","0101","0010","0100","0110","0010","0011","0101","0011","0011","0110","0101","0010","0010","0011","0011","0010","0010","0011","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0100","0011","0100","0110","0110","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0010","0011","0011","0101","0111","1001","1010","1001","1000","0110","0110","0110","0110","0101","0001","0000","0000","0001","0010","0011","0100","0011","0011","0011","0010","0100","0110","0101","0100","0011","0011","0100","0101","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0111","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","1000","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0111","0111","0111","0110","0111","0110","0111","0110","0110","1000","0111","0111","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0101","0101","0101","0101","0100","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0001","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0000","0000","0001","0000","0000","0000"),
("0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0100","0011","0110","0111","0111","0110","0101","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0100","0010","0100","0101","0011","0011","0101","0011","0011","0101","0011","0100","0110","0110","0011","0101","0111","0100","0100","1000","0110","0011","0100","0011","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0101","0111","0011","0110","1001","0101","0101","1001","0111","0100","1000","0101","0011","0110","0111","0011","0101","1000","0011","0100","1000","0100","0011","0111","0110","0010","0110","0111","0011","0111","1001","0101","0010","0011","0010","0010","0010","0010","0100","0100","0100","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0100","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0111","0111","0110","0100","0011","0011","0011","0011","0011","0010","0011","0101","0100","0101","0110","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0101","0101","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0111","0111","0110","0111","0111","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0110","1000","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0110","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0101","0101","0101","0101","0110","0100","0011","0010","0010","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0010","0100","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","0011","0010","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0001","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0001","0010","0011","0011","0011","0011"),
("0110","0111","0111","0111","0111","0111","0110","0111","0111","0111","0100","0011","0110","0111","0111","0110","0011","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0011","0100","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","1000","0111","0011","0111","1000","0100","0110","0111","0010","0100","0111","0101","0011","0111","0101","0011","0111","0111","0011","0101","1000","0011","0100","1000","0101","0100","1001","0111","0010","0011","0010","0011","0010","0010","0011","0100","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0100","0011","0100","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0010","0010","0010","0010","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0101","0110","0101","0101","0110","0101","0101","0110","0110","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0101","0110","0101","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0101","0110","0110","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","1000","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0111","1000","0111","0111","1000","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0101","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0100","0100","0101","0110","0110","0101","0100","0011","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0100","0100","0011","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0010","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0011","0011","0100","0100","0100"),
("0100","0011","0011","0100","0100","0100","0011","0100","0100","0101","0100","0011","0101","0101","0101","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0011","0011","0011","0100","0100","0011","0100","0100","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0011","0100","0010","0011","0100","0011","0011","0100","0011","0010","0100","0100","0010","0011","0100","0010","0100","0101","0011","0010","0011","0010","0010","0010","0011","0100","0100","0101","0100","0101","0101","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0100","0011","0011","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0011","0100","0101","0101","0101","0110","0110","0110","0110","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0110","0101","0110","0110","0101","0110","0110","0110","0110","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0110","0110","0110","0111","0110","0111","0111","0110","0111","0110","0110","0110","0101","0110","0110","0110","0111","0110","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0111","0110","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0100","0101","0101","0110","0110","0110","0101","0100","0011","0011","0011","0010","0001","0001","0010","0001","0001","0010","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0011","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0001","0011","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0100","0100","0100","0100"),
("0100","0001","0011","0010","0010","0001","0000","0001","0010","0100","0011","0010","0011","0011","0100","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0001","0010","0010","0011","0011","0010","0001","0001","0011","0011","0011","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0100","0011","0101","0101","0101","0101","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0100","0011","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0101","0101","0110","0101","0110","0110","0110","0111","0110","0110","0110","0110","0111","0110","0111","0111","0110","0111","0111","0110","0111","0110","0111","0110","0110","1000","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0110","0111","0101","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0100","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0010","0010","0010","0010","0001","0001","0010","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0000","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0000","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0010","0011","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0101","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0100","0100","0011","0100"),
("0100","0001","0010","0010","0010","0001","0001","0001","0010","0011","0011","0010","0010","0100","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0000","0000","0010","0111","1000","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0101","0100","0100","0101","0100","0100","0101","0100","0100","0100","0101","0100","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0100","0100","0011","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0101","0100","0101","0100","0100","0101","0101","0101","0100","0100","0100","0101","0100","0101","0100","0101","0100","0100","0101","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0101","0100","0101","0100","0100","0101","0101","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0110","0110","0101","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0110","0111","0111","0111","0111","0110","0111","0110","0110","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0100","0100","0101","0101","0101","0101","0101","0011","0011","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0000","0000","0001","0001","0010","0010","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0010","0010","0001","0010","0010","0010","0001","0010","0010","0001","0010","0010","0010","0001","0010","0010","0001","0001","0010","0010","0011","0011","0011","0011","0100"),
("0100","0001","0010","0001","0010","0001","0001","0001","0001","0010","0010","0010","0010","0101","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0001","0000","0001","0001","0000","0000","0010","0111","1000","0011","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0101","0101","0011","0110","0110","0101","0110","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0100","0101","0101","0101","0011","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0101","0111","0111","0110","0111","0111","0111","1000","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","1000","0111","0110","0111","0110","0111","0111","0110","0111","0110","0111","0111","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0100","0100","0101","0101","0100","0101","0101","0011","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0010","0001","0000","0000","0000","0001","0011","0010","0011","0011","0011","0011","0011","0100","0011","0100","0100","0100","0100","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0011","0010","0011","0011","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0011","0010","0010","0011","0011","0001","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0011","0010","0010","0011","0011","0100","0011"),
("0100","0001","0010","0001","0010","0001","0001","0001","0010","0010","0010","0001","0100","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0101","0101","0101","0110","0110","0100","0011","0011","0011","0100","0101","0100","0010","0010","0010","0010","0010","0001","0010","0111","1000","0011","0010","0010","0010","0011","0011","0010","0010","0010","0001","0011","0110","0100","0010","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0101","0101","0100","0100","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0011","0011","0100","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0011","0011","0101","0101","0101","0101","0101","1000","0110","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0011","0100","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0101","0100","0100","0100","0100","0101","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0101","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0110","0101","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0111","0111","0111","0111","0110","0111","0110","0111","1000","0110","0111","0110","0110","0111","0110","0111","0111","0110","0111","0110","0011","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0100","0100","0100","0101","0101","0101","0101","0100","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0001","0000","0000","0000","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0100","0011","0011","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0001","0001","0001","0010","0001","0000","0001","0010","0001","0001","0010","0010","0001","0010","0010","0001","0010","0011","0010","0010","0010","0010","0011","0010","0000"),
("0101","0001","0010","0010","0010","0001","0001","0001","0010","0011","0010","0010","0101","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0111","0111","1000","1000","1000","1000","0101","0110","1001","1001","1001","1001","1000","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0001","0010","0101","0100","0011","0011","0100","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0001","0101","0110","0101","0101","0110","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0101","0101","0101","0100","0100","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0110","0101","0100","0101","0111","1000","0111","0110","0111","0111","0110","0111","0110","0111","1000","0110","0111","0110","0110","0111","0111","0111","0111","0110","0111","0110","0111","1000","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0100","0011","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0100","0100","0101","0101","0101","0101","0110","0100","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0010","0010","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0100","0011","0100","0100","0011","0011","0011","0011","0100","0100","0100","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0010","0010","0010","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0101","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0100","0011","0000"),
("0101","0010","0010","0010","0010","0001","0001","0001","0010","0100","0010","0011","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0111","1000","1001","1001","1001","1001","1010","1010","1010","1010","1010","0111","0110","1001","1001","1001","1000","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0001","0101","0101","0011","0011","0100","0011","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0001","0011","0101","0110","1000","0110","0101","0101","0101","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0100","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0100","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0110","0101","0101","0101","0110","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","1000","0110","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0110","0110","0111","0110","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0101","0100","0101","0110","0101","0101","0110","0101","0101","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0000","0001","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0011","0011","0011","0100","0100","0100","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0010","0001","0010","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0101","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0001","0011","0011","0011","0010","0001"),
("0101","0011","0011","0010","0010","0001","0001","0001","0010","0010","0010","0101","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0000","0011","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1001","1010","1001","1010","1001","1001","1001","0110","1000","1010","1010","1000","0101","1001","1010","0111","0101","0011","0100","0100","0100","0100","0100","0011","0011","0100","0011","0100","0100","0100","0011","0100","0011","0010","0010","0100","0101","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0100","0011","0011","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0011","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0001","0110","0111","0110","0101","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0110","0101","0101","0101","0101","0110","0110","0111","0111","0110","0111","0111","0111","0111","0110","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0111","0110","0110","0111","0111","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0101","0110","0110","0101","0100","0100","0100","0100","0110","0101","0101","0110","0101","0101","0101","0101","0101","0101","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0001","0000","0010","0010","0011","0100","0011","0011","0101","0110","0101","0011","0100","0100","0100","0100","0011","0100","0101","0100","0011","0100","0100","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0101","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0001","0010","0010","0010","0010","0001"),
("0100","0100","0100","0100","0011","0010","0010","0011","0011","0011","0100","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0001","0011","1000","1001","0110","0010","0110","1001","0111","0011","0110","1001","0111","0100","0111","1000","1000","1010","0111","0101","1010","0101","0111","1010","0100","1000","1010","1010","1001","0101","1001","1000","0100","0011","0011","0100","0100","0100","0100","0100","0110","0110","0011","0010","0100","0100","0100","0100","0011","0011","0001","0100","0101","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0010","0010","0010","0011","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0100","0101","0100","0101","0100","0100","0100","0100","0101","0101","0101","0101","0100","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0110","0110","0101","0101","0101","0101","0101","0111","0111","0111","0111","0110","0111","0111","0111","1000","0111","0111","0111","0110","0111","0110","0110","0111","0110","0111","0111","0110","0110","0100","0110","0111","0110","0011","0001","0001","0011","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0010","0001","0010","0010","0001","0011","0101","0101","0101","0110","0110","0110","0101","0101","0101","0101","0101","0100","0100","0100","0100","0010","0001","0001","0001","0001","0001","0000","0001","0000","0000","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0000","0001","0011","0010","0100","0100","0011","0011","1000","1001","0110","0011","0100","0100","0100","0011","0011","1000","1001","0111","0100","1010","1011","0111","0011","0100","0100","0011","0011","0011","0011","0011","0011","0101","0110","0101","0011","0101","0110","0100","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0101","0010","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0001","0010","0010","0010","0010","0000"),
("0011","0100","0010","0010","0010","0010","0010","0010","0010","0011","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0010","0010","0100","1000","1001","0101","0000","0110","1001","0110","0000","0101","1001","0111","0000","0101","1001","1000","1001","0110","0101","1010","0110","0111","1010","0111","1001","1010","1010","1001","0110","0110","0100","0011","0011","0011","0100","0100","0100","0011","0110","1001","0110","0010","0011","0100","0100","0011","0011","0011","0011","0100","0101","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0011","0011","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0011","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0101","0101","0101","0100","0100","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0111","0111","0111","0111","0111","1000","0111","0111","1000","0111","0111","1000","0111","1000","0111","0110","0110","0110","0100","0011","0101","0110","0110","0100","0011","0011","0100","0100","0100","0100","0100","0101","0101","0101","0100","0101","0101","0100","0010","0001","0001","0010","0011","0100","0101","0101","0101","0101","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0011","0010","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0000","0010","0010","0011","0100","0100","0011","0101","1001","1000","0100","0011","0100","0100","0100","0011","0101","1001","1000","0100","0111","1100","1011","0101","0011","0100","0011","0011","0011","0011","0011","0011","0100","1000","1000","0110","0100","1001","1001","0110","0011","0100","0011","0011","0011","0011","0011","0011","0011","0111","1000","0110","0010","0011","0011","0100","0111","0110","0011","0010","0001","0001","0001","0010","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0001","0010","0010","0001","0010","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0101","0010","0010","0001","0001","0010","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0001","0010","0010","0010","0010","0000"),
("0101","0101","0010","0010","0010","0010","0001","0001","0001","0100","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0010","0010","0100","1001","1000","1000","0110","1000","1001","1000","0110","0111","1001","1000","0101","0111","1001","1001","1001","1000","0111","1010","1001","1001","1010","1010","1001","1001","1001","1001","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0100","0110","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0100","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0101","0101","0101","0100","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0100","0101","0110","0101","0101","0101","0101","0101","0101","0101","0110","0111","0110","0110","0111","0110","0110","0110","0101","0101","0110","0101","0110","0110","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0011","0100","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0010","0000","0001","0010","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0011","0010","0100","0100","0011","0010","0101","0110","0101","0011","0100","0100","0100","0100","0011","0111","1001","1000","0011","1001","1100","1001","0011","0100","0100","0011","0011","0011","0011","0011","0011","0110","1001","1000","0100","0111","1001","1000","0100","0011","0011","0011","0011","0011","0011","0011","0011","0101","1001","1000","0100","0011","0100","0011","0111","1000","0111","0011","0010","0000","0001","0010","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0110","0111","0101","0001","0010","0010","0001","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0101","0010","0010","0001","0001","0010","0001","0001","0010","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0001","0010","0010","0010","0010","0000"),
("0110","0101","0010","0010","0010","0010","0010","0000","0001","0100","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0010","0010","0100","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1010","1010","1010","1010","1010","1001","1000","1000","0101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0100","0101","0100","0101","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0100","0100","0100","0101","0101","0100","0100","0100","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0101","0100","0100","0101","0100","0101","0101","0100","0101","0101","0101","0100","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0101","0100","0101","0100","0011","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0100","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0100","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0011","0100","0110","0110","0110","0110","0110","0101","0100","0100","0011","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0100","0010","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0010","0010","0011","0100","0100","0011","0010","0010","0010","0010","0011","0100","0100","0100","0011","0100","1001","1001","0110","0101","1011","1011","0110","0011","0100","0100","0011","0011","0011","0011","0100","0011","1000","1000","0111","0011","1001","1001","0111","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","1001","0111","0011","0011","0011","0011","1000","1000","0101","0011","0010","0001","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","1000","0111","0100","0001","0010","0010","0010","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0101","0010","0010","0001","0001","0010","0001","0010","0010","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0001","0010","0010","0010","0010","0000"),
("0110","0101","0010","0001","0010","0010","0010","0000","0011","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0011","0011","0011","0011","0011","0100","0100","0011","0010","0010","0100","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1010","1010","1010","1010","1001","1010","1001","1001","1000","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0100","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0100","0101","0101","0100","0100","0100","0100","0101","0100","0100","0100","0101","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0100","0011","0010","0101","0101","0110","0100","0100","0101","0101","0101","0101","0101","0011","0011","0011","0011","0011","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0011","0011","0010","0010","0010","0011","0010","0010","0010","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0100","0011","0010","0100","0010","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0011","0011","0011","0101","0101","0011","0100","1000","1000","0100","0011","0100","0011","0011","0011","0011","0011","0011","0100","1000","1000","0101","0101","1001","1000","0101","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0101","1000","1000","0100","0011","0011","0010","0001","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0101","0111","0110","0011","0010","0010","0010","0010","0101","0110","0110","0110","0110","0110","0110","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0101","0100","0010","0001","0001","0001","0001","0001","0010","0010","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0001","0010","0011","0010","0010","0001"),
("0110","0101","0011","0011","0011","0100","0100","0011","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0001","0011","0010","0010","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","1000","1001","0111","0100","0111","1001","1000","0110","0111","1001","1000","0110","0111","1001","1001","1001","1000","0110","1001","0111","0110","1001","1001","1000","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0100","0100","0011","0011","0011","0100","0100","0101","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0101","0101","0100","0100","0100","0101","0100","0100","0101","0100","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0110","0110","0100","0100","0011","0011","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0010","0000","0000","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0011","0010","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0110","0111","0110","0010","0011","0000","0000","0001","0011","0011","0011","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0110","0110","0110","0110","0110","0110","0101","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0010","0001","0001"),
("0101","0100","0100","0101","0101","0101","0101","0100","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0001","0001","0001","0001","0010","0011","0011","0011","0100","0011","0100","0011","0010","0010","0100","1000","1001","0110","0000","0101","1001","0111","0000","0101","1001","0111","0000","0101","1001","1001","1001","0111","0100","1001","0110","0101","1001","1000","0100","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0100","0011","0011","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0100","0100","0101","0100","0101","0101","0100","0100","0101","0101","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0101","0101","0100","0011","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0101","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0100","0100","0011","0010","0011","0111","1000","1000","0100","0011","0101","0101","0100","0100","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0100","0100","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0010","0001","0001","0001","0001","0001","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0010","0011","0100","0011","0011","0100","0011","0100","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","0011","0011","0001","0001","0010","0001","0001","0001","0001","0001","0010","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0100","0110","0110","0110","0110","0110","0110","0100","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0000","0000","0000","0000","0001","0001","0010","0010","0010","0010"),
("0110","0110","0110","0110","0110","0110","0101","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0010","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","1000","1001","0111","0101","0111","1001","0111","0100","0110","1001","0111","0011","0110","1001","1000","1000","0111","0101","1001","1000","1000","1000","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0100","0101","0100","0100","0100","0011","0011","0010","0011","0100","0101","0101","0100","0100","0011","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0100","0101","0100","0100","1001","1100","1100","0101","0010","0110","1100","1100","1011","0011","0100","0101","0100","0100","0011","0111","1001","1001","0011","0010","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0101","0100","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0101","0100","0101","0100","0100","0100","0100","0101","0100","0101","0101","0101","0100","0101","0101","0100","0100","0100","0100","0100","0101","0100","0100","0100","0101","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0101","0101","0101","0101","0100","0101","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0101","0100","0101","0101","0100","0100","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0011","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0010","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0000","0001","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0001","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0001","0010","0101","0110","0110","0110","0110","0101","0101","0010","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0000","0000","0000","0001","0001","0010","0001","0010","0100"),
("0110","0110","0110","0110","0110","0101","0100","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1000","1000","1000","1000","1001","1001","1000","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0010","0001","0010","0010","0010","0010","0011","0011","0011","0100","0101","0101","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0100","0101","0101","0100","0100","0011","0010","0010","0010","0011","0100","0101","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","1000","1100","1101","1001","0010","0100","1010","1100","1100","0110","0011","0101","0101","0100","0100","0110","1011","1011","1001","0010","0100","0100","0101","0100","0100","0100","0100","0101","0101","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0100","0101","0110","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0101","0100","0100","0100","0100","0011","0010","0011","0101","0101","0011","0001","0000","0001","0001","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0010","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0000","0000","0001","0001","0001","0011","0100","0011","0100","0011","0100","0011","0100","0011","0100","0100","0100","0011","0100","0011","0011","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0001","0011","0110","0110","0110","0110","0110","0101","0101","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0010","0010"),
("0110","0110","0110","0110","0101","0101","0011","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1000","1000","1000","1001","0111","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0001","0001","0001","0010","0010","0001","0010","0010","0001","0010","0010","0011","0010","0010","0001","0010","0011","0010","0010","0010","0011","0100","0100","0100","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0100","0110","0111","0111","0111","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0110","1100","1100","1011","0011","0010","0111","1100","1100","1010","0010","0100","0101","0100","0100","0101","1011","1011","1010","0100","0011","0101","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0110","0111","0111","0100","0010","0011","0100","0100","0100","0010","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0100","0101","0101","0101","0101","0100","0100","0100","0101","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0101","0100","0101","0100","0100","0101","0101","0100","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0011","0011","0011","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0100","0010","0010","0011","0011","0100","0011","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0101","0100","0100","0100","0101","0100","0100","0100","0010","0011","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0100","0101","0101","0010","0001","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0010","0001","0000","0001","0000","0001","0000","0000","0000","0001","0001","0000","0001","0001","0001","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0100","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0100","0110","0110","0110","0101","0101","0101","0011","0000","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0010","0001"),
("0110","0110","0110","0110","0101","0100","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","0111","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0001","0010","0011","0010","0010","0011","0010","0010","0001","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0001","0010","0011","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0101","0111","0111","0111","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0101","0111","0111","0101","0001","0011","1001","1011","1011","0101","0011","0101","0101","0101","0100","1000","1010","1010","0110","0001","0100","0101","0101","0100","0101","0100","0100","0101","0100","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","1101","1110","1101","0101","0010","0110","0101","1001","0111","0010","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","1010","1001","1000","0010","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0011","0001","0000","0001","0001","0011","0100","0100","0100","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0011","0011","0011","0011","0011","0101","0100","0100","0101","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0101","0101","0011","0001","0001","0001","0011","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0001","0010","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0100","0011","0011","0011","0011","0011","0010","0100","0100","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0111","1000","0101","0001","0000","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0011","0100","0100","0100","0100","0100","0010","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0100","0100","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0100","0101","0110","0110","0101","0101","0101","0101","0010","0000","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0001","0001","0001"),
("0110","0110","0110","0110","0101","0011","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0001","0001","0010","0111","1000","1000","0110","0010","0010","0011","0011","0011","0011","0011","0100","0101","0100","0100","0110","0110","0101","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0011","0011","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0001","0000","0010","0100","0101","0101","0101","0101","0100","0100","0011","0100","0101","0101","0101","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0100","0100","0011","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0001","0001","0001","0001","0011","0010","0011","0011","0011","0010","0100","0101","0101","0101","0010","0010","0010","0011","0001","0011","0101","0101","0101","0100","0100","0101","0100","0101","0101","0100","0100","0101","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","1001","1101","1110","1010","0010","0100","1001","0101","1000","0100","0011","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","1010","1101","1101","0111","0010","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0001","0001","0010","0010","0100","0100","0101","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0011","0010","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0011","0101","0101","0100","0101","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0010","0001","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0001","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0011","0001","0000","0001","0010","0010","0001","0010","0011","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0111","1000","0100","0000","0010","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0010","0001","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0000","0001","0010","0001","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0011","0010","0001","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0101","0101","0110","0110","0101","0101","0101","0100","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0000","0001","0001","0001"),
("0110","0110","0101","0101","0100","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0000","0000","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0111","1000","1000","0110","0001","0000","0000","0001","0001","0000","0000","0110","0111","0111","0111","0101","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0010","0001","0001","0010","0010","0001","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0010","0001","0010","0010","0010","0001","0010","0010","0001","0001","0010","0001","0010","0010","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0001","0001","0010","0010","0100","0011","0011","0011","0100","0011","0001","0010","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0011","0011","0011","0011","0011","0100","0100","0101","0101","0100","0100","0101","0101","0100","0101","0100","0100","0100","0100","0100","0101","0100","0101","0101","0101","0101","0100","0101","1100","1101","1101","0101","0011","0111","1001","0101","0110","0010","0100","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0110","1100","1100","1011","0011","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0001","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","1010","1010","1010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0101","0100","0011","0100","1010","1010","1001","0011","0011","0101","0101","0101","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0010","0010","0010","0100","0100","0011","0100","0011","0010","0010","0010","0011","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0010","0010","0010","0011","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0001","0001","0010","0010","0010","0011","0010","0100","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0101","0111","0111","0101","0001","0011","0100","0100","0100","0100","0100","0100","0011","0010","0011","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0010","0011","0010","0001","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0001","0010","0100","0101","0100","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0110","0101","0110","0110","0101","0101","0101","0011","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0010","0010","0001","0001","0010","0001","0001","0001","0001"),
("0110","0110","0101","0100","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0001","0000","0000","0001","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0111","1000","1000","0110","0001","0000","0000","0001","0001","0000","0001","0110","0111","1000","0111","0011","0001","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0001","0001","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0001","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0100","0101","0101","0101","0101","0101","0101","0100","0100","0101","0100","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","1001","1101","1101","1010","0011","0100","1010","1000","0010","0010","0011","0101","0100","0101","0100","0011","0100","0101","0101","0100","0100","0100","0101","0100","0101","0100","0100","1010","1100","1100","0111","0010","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0001","0001","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0100","0011","0111","1010","1010","0111","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","1000","1100","1100","1001","0010","0100","0100","0100","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0100","0100","0011","0001","0100","0100","0100","0011","0011","0010","0010","0011","0011","0100","0100","0100","0100","0100","0101","0101","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0011","0100","0101","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0010","0001","0010","0010","0010","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0110","0111","0111","0101","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0011","0010","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0010","0100","0010","0001","0010","0001","0000","0000","0001","0000","0001","0001","0000","0001","0000","0000","0000","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0001","0000","0001","0010","0011","0101","0110","1000","1000","1000","0111","0111","0110","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","0100","0110","0101","0101","0101","0101","0001","0000","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0010","0010","0010"),
("0110","0110","0101","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0010","0010","0011","0010","0000","0000","0000","0000","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","0111","0111","0110","0001","0000","0000","0001","0010","0000","0001","0110","1000","0111","0100","0010","0001","0010","0010","0010","0010","0011","0010","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0001","0001","0010","0010","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0001","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0011","0101","0110","0110","0100","0011","0011","0111","0101","0011","0011","0100","0101","0100","0100","0011","0010","0011","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","1010","1010","1010","0011","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0010","0001","0000","0000","0000","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0101","1010","1010","1001","0100","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","1011","1100","1100","0101","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0100","0101","0101","0101","0100","0100","0100","0011","0111","1010","1010","0110","0010","0100","0100","0100","0100","0011","0010","0010","0011","0010","0011","0100","0100","0100","0100","0011","0101","0101","0011","0100","0101","0100","0100","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0010","0011","0010","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0110","0111","0111","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0010","0100","0010","0010","0011","0010","0000","0001","0000","0000","0000","0000","0000","0001","0000","0000","0000","0010","0011","0011","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0100","0100","0011","0010","0110","0111","1000","0111","0111","0111","1000","0101","0100","0111","1000","0111","0110","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0010","0100","0110","0101","0101","0101","0100","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0010","0001","0001"),
("0101","0101","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0101","0101","0101","0101","0100","0010","0101","0101","0100","0001","0010","0011","0011","0010","0011","0010","0000","0000","0000","0000","0000","0000","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","1000","0111","0110","0001","0001","0000","0010","0011","0001","0001","0110","0110","0110","0101","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0001","0001","0010","0001","0001","0000","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0001","0010","0010","0010","0001","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0011","0100","0011","0010","0100","0100","0101","0101","0100","0100","0011","0011","0010","0010","0010","0011","0100","0101","0101","0101","0101","0101","0100","0001","0010","0010","0010","0011","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0011","0001","0001","0000","0000","0001","0011","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0101","0100","0011","0101","1000","1000","0110","0001","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0101","0101","0100","0100","0100","0011","1000","1100","1100","1010","0010","0100","0101","0101","0101","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0110","1011","1010","1001","0011","0011","0100","0100","0100","0011","0011","0010","0010","0010","0011","0011","0100","0100","0101","0100","0101","1100","1011","0011","0011","0101","0100","1010","1100","0110","0011","0100","0100","0100","0011","0011","0010","0001","0011","0010","0010","0101","0101","0100","1000","1000","0011","0011","0100","0011","0100","0011","0010","0001","0010","0011","0010","0100","0011","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0100","0100","0100","0100","0011","0010","0010","0001","0001","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0010","0100","0010","0010","0100","0011","0000","0001","0000","0001","0010","0010","0001","0001","0000","0000","0000","0010","0100","0100","0001","0000","0000","0000","0010","0010","0001","0100","0111","1000","1000","0111","0111","0111","0110","0110","0110","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0110","0110","0101","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0110","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0001","0001","0010","0100","0110","0101","0101","0101","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0100","0100","0011","0010","0101","0101","0011","0001","0011","0011","0001","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","0111","0111","0110","0001","0001","0000","0001","0010","0001","0001","0110","0111","0110","0111","0110","0100","0101","0100","0011","0100","0101","0100","0011","0101","0100","0100","0100","0100","0011","0011","0011","0011","0010","0011","0010","0001","0010","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0100","0011","0011","0010","0010","0010","0010","0100","0011","0011","0010","0001","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0001","0001","0011","0011","0010","0010","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0010","0011","0100","0100","0101","0101","0100","0100","0101","0101","0101","0100","0100","0101","0101","0101","0101","0100","0010","0001","0001","0001","0001","0010","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0101","0100","0100","0100","0100","0010","0011","0100","0100","0011","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","1001","1010","1010","0110","0001","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","1001","1101","1001","0010","0100","0100","0110","1100","1100","0100","0100","0100","0100","0100","0100","0100","0010","0101","0100","0010","0011","0100","0100","0111","1101","1011","0011","0100","0100","0100","0100","0011","0010","0010","0010","0010","0100","0100","0011","0011","0100","0101","0101","0101","0101","0101","0101","0110","0101","0101","0100","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0100","0100","0100","0011","0010","0011","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0100","0010","0010","0100","0011","0000","0001","0000","0001","0010","0010","0010","0001","0000","0000","0000","0010","0100","0011","0010","0010","0011","0101","0110","0101","0100","0111","0111","0111","0110","0100","0110","0111","1000","1000","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","1000","1000","1000","0111","0111","0110","0101","0101","0101","0100","0100","0011","0011","0011","0110","0011","0010","0001","0000","0000","0000","0000","0001","0000","0000","0000","0001","0010","0010","0010","0010","0010","0100","0101","0101","0101","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0001","0001","0001","0010"),
("0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","0111","0111","0110","0001","0000","0000","0001","0001","0000","0001","0101","1000","0110","0110","0111","0111","0101","0100","0011","0100","0011","0011","0011","0100","0011","0100","0010","0011","0100","0100","0110","0101","0100","0100","0100","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0100","0011","0011","0100","0011","0011","0011","0011","0010","0010","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0100","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0011","0010","0001","0000","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0001","0001","0001","0010","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0100","0100","0100","0010","0011","0011","0011","0001","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","1011","1100","0101","0011","0101","0100","1001","1101","1001","0011","0101","0100","0101","0100","0100","0011","0100","1001","0100","0010","0100","0101","0100","1010","1101","0111","0010","0100","0100","0100","0100","0011","0010","0010","0010","0011","0100","0100","0011","0011","0101","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0011","0010","0010","0010","0011","0010","0010","0001","0000","0000","0001","0001","0001","0000","0000","0010","0100","0010","0010","0101","0011","0000","0001","0000","0001","0001","0001","0010","0001","0000","0000","0001","0010","0100","0110","0111","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","1000","0111","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","0111","0111","0110","0101","0100","0100","0010","0010","0101","0011","0010","0001","0000","0000","0000","0000","0001","0000","0000","0000","0001","0011","0011","0010","0010","0010","0100","0110","0101","0101","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","0111","0111","0110","0001","0001","0001","0001","0011","0001","0001","0100","0110","0111","0110","0110","0110","0101","0110","0111","0110","0111","0110","0100","0101","0100","0101","0101","0011","0011","0100","0101","0101","0101","0101","0101","0011","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0000","0000","0001","0001","0001","0001","0000","0000","0001","0001","0000","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0100","0100","0011","0100","0011","0011","0100","0011","0011","0011","0010","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0101","0111","0101","0011","0011","0010","0010","0010","0011","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0101","0100","0100","0100","0100","0011","0010","0010","0011","0010","0010","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0001","0001","0001","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0011","0010","0100","0100","0010","0100","0100","0010","0101","0110","0011","0100","0101","0101","0101","0100","0100","0001","0010","0011","0100","0100","0100","0100","0100","1010","1010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0101","0101","0110","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0001","0001","0000","0000","0000","0000","0010","0100","0011","0010","0100","0011","0000","0001","0000","0000","0001","0001","0010","0010","0011","0101","0110","0111","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","1000","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0110","0101","0100","0101","0100","0011","0001","0000","0000","0000","0001","0001","0001","0000","0000","0001","0011","0011","0010","0011","0010","0100","0110","0101","0101","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","1000","0111","0110","0001","0001","0001","0001","0010","0000","0001","0100","0110","0111","0110","0110","0110","0100","0101","0100","0011","0101","0100","0011","0100","0100","0100","0100","0010","0010","0011","0100","0011","0011","0101","0100","0010","0010","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0010","0001","0010","0001","0010","0010","0010","0010","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0011","0100","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0011","0010","0010","0011","0100","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0100","1000","0110","0011","0010","0100","1010","1011","1000","0100","0011","0011","0011","0010","0010","0010","0011","0100","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0101","0100","0101","0101","0101","0101","0100","0101","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0011","0100","0011","0011","0011","0010","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0101","0101","0101","0100","0101","0100","0100","0100","0100","0100","0100","0101","0100","0101","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0011","0011","0100","0100","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0010","0010","0100","0101","0101","0100","0011","0010","0010","0010","0010","0100","0100","0100","0101","0101","0100","0100","0011","0011","0100","0100","0100","0100","0100","0101","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0010","0001","0010","0000","0000","0001","0100","0011","0010","0100","0011","0000","0001","0001","0010","0010","0001","0010","0110","0111","1000","1000","1000","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","1000","0111","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0111","0111","0110","0101","0100","0010","0000","0000","0001","0001","0000","0000","0001","0011","0011","0011","0011","0010","0100","0101","0101","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0011","0010","0001","0001","0010","0010","0001","0001","0001","0001","0010","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0010","0001","0001"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0111","1000","0111","0110","0001","0001","0001","0000","0001","0000","0001","0110","0110","0111","0110","0101","0101","0110","0101","0001","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0100","0011","0100","0011","0100","0100","0001","0010","0001","0000","0001","0010","0010","0011","0010","0010","0010","0011","0011","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010","0010","0001","0010","0010","0010","0010","0011","0011","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0101","0110","0111","0110","0110","0111","0111","1000","1000","0111","0111","0111","0100","0010","0010","0010","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0101","0100","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0001","0001","0011","0010","0010","0001","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0101","0110","0100","0011","0011","0011","1000","1011","1001","0101","0011","0011","0110","1011","1010","0111","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0011","0011","0011","0011","0010","0010","0010","0010","0011","0100","0011","0100","0100","0011","0100","0011","0011","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0100","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0011","0100","0100","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0011","0010","0011","0010","0000","0001","0010","0010","0010","0100","0101","0100","0110","0111","0111","0110","0101","0101","0110","0110","0111","0111","0111","0101","0100","0110","0111","1000","0111","0111","1000","1000","1000","0111","0111","1000","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0100","0011","0010","0001","0000","0000","0001","0000","0000","0001","0011","0100","0011","0011","0011","0100","0101","0101","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0110","0111","0111","0111","0010","0001","0001","0001","0001","0001","0001","0101","0110","0100","0101","0100","0100","0101","0100","0010","0000","0001","0000","0000","0000","0000","0001","0000","0000","0001","0101","0100","0011","0100","0010","0010","0010","0010","0001","0001","0010","0100","0101","0011","0010","0001","0010","0011","0010","0010","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0011","0011","0010","0011","0011","0011","0101","0100","0110","0110","0110","0110","0111","0111","0111","0101","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0011","0011","0100","0011","0010","0011","0100","0011","0011","0011","0011","0011","0011","0010","0100","1010","1011","0111","0011","0011","0010","0100","1001","1011","1000","0100","0010","0011","1000","1011","1001","0100","0011","0011","0011","0010","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0100","0100","0011","0011","0010","0010","0011","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0011","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0101","0101","0101","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0101","0100","0101","0101","0100","0101","0101","0100","0100","0100","0100","0100","0011","0010","0011","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0001","0000","0011","0100","0111","1001","1001","1000","1000","0111","0111","0110","0110","0110","0110","0111","0111","0111","1000","0111","0111","0111","0111","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","1000","1000","0111","1000","0111","0111","0111","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0100","0011","0011","0010","0001","0001","0000","0000","0000","0001","0000","0000","0001","0010","0100","0011","0011","0010","0100","0101","0101","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0010","0001","0001","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0110","0111","0111","0111","0010","0001","0001","0001","0001","0001","0001","0011","0101","0100","0100","0111","0100","0011","0011","0010","0000","0001","0000","0000","0000","0000","0000","0000","0000","0001","0100","0101","0011","0100","0010","0011","0011","0100","0010","0010","0100","0101","0101","0100","0011","0001","0010","0010","0010","0010","0001","0001","0010","0011","0010","0001","0010","0010","0010","0001","0001","0001","0010","0010","0001","0011","0101","0011","0010","0010","0001","0001","0001","0001","0001","0001","0011","0011","0011","0011","0101","0101","0100","0100","0110","0111","0111","1000","0111","0101","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0010","0010","0001","0010","0001","0001","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0011","0010","0011","0010","0010","0010","0011","0011","0011","0010","0011","0011","0100","0011","0010","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0111","1011","1010","0110","0011","0011","0011","0110","1010","1010","0101","0011","0010","0100","0100","0011","0010","0001","0001","0010","0010","0010","0011","0011","0010","0001","0001","0001","0011","0100","0100","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0010","0011","0011","0010","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0010","0010","0001","0001","0001","0010","0011","0011","0011","0010","0010","0010","0011","0010","0010","0011","0011","0011","0010","0100","0100","0011","0101","0110","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0111","1000","1000","0110","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0100","0011","0010","0010","0010","0011","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0010","0100","0011","0011","0011","0100","0101","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0001","0101","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0110","0111","1000","0111","0010","0001","0001","0001","0001","0001","0001","0011","0110","0101","0011","0101","0100","0010","0101","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0100","0100","0100","0100","0001","0100","0011","0100","0010","0010","0011","0100","0100","0100","0011","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0001","0001","0001","0010","0010","0001","0010","0100","0010","0001","0001","0001","0001","0001","0001","0001","0010","0011","0010","0100","0011","0011","0011","0011","0100","0110","1000","1001","1000","0100","0010","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0001","0001","0010","0010","0011","0010","0010","0010","0001","0001","0001","0001","0001","1000","1000","0100","0011","0010","0001","0001","0001","0010","0011","0011","0011","0011","0011","0100","1001","1011","1000","0100","0011","0011","0011","0100","0011","0010","0001","0001","0001","0011","0100","0011","0010","0010","0010","0010","0001","0000","0001","0001","0000","0001","0011","0100","0110","0110","0110","0110","0110","0110","0011","0001","0001","0001","0001","0001","0010","0101","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0101","0101","0101","0101","0100","0101","0100","0100","0101","0100","0100","0101","0101","0101","0100","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0101","0100","0101","0100","0101","0101","0101","0100","0100","0100","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0001","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0101","0110","0111","0111","0111","0111","0111","0111","0111","1000","0111","0100","0111","0111","0111","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","1000","0111","0111","0111","0110","0110","0101","0100","0100","0011","0011","0010","0001","0001","0001","0010","0010","0001","0001","0000","0001","0001","0001","0000","0001","0000","0000","0000","0001","0100","0011","0011","0011","0101","0101","0011","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0010","0001","0001","0010","0011","0011","0011","0010","0001","0001","0010","0010","0010","0001","0101","0111","0110","0110","0111","0110","0110","0110","0111","0110","0110","0110","0110","0111","0111","0111","0110","0111","0110"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0110","0110","1000","0111","0010","0001","0001","0001","0001","0001","0001","0100","0110","0110","0011","0011","0100","0100","0100","0011","0001","0001","0000","0000","0000","0000","0000","0000","0000","0010","0100","0011","0100","0010","0001","0011","0010","0100","0011","0001","0010","0011","0010","0010","0011","0010","0001","0011","0001","0000","0010","0011","0001","0001","0001","0010","0010","0001","0010","0000","0001","0001","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0011","0011","0100","0100","0010","0001","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0110","0110","0011","0010","0001","0001","0010","0010","0010","0011","0100","0011","0011","0011","0010","0101","0110","0100","0010","0001","0001","0001","0011","0011","0011","0010","0010","0010","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0001","0010","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0011","0010","0010","0010","0010","0010","0011","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0100","0011","0011","0011","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0100","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0010","0010","0011","0010","0001","0001","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0011","0010","0010","0011","0011","0011","0100","0100","0110","0111","0111","1000","1000","0111","0100","0011","0101","0111","1000","0111","1000","1000","0111","0111","1000","1000","0111","1000","1000","1000","0111","1000","0111","0111","1000","1000","0111","0111","0111","0111","0110","0110","0110","0101","0100","0011","0010","0010","0001","0001","0001","0000","0000","0001","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0010","0001","0100","0101","0010","0010","0011","0011","0011","0011","0100","0011","0011","0010","0010","0001","0010","0101","0110","0111","0111","0110","0101","0011","0010","0010","0010","0010","0001","0101","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0101","0111","0111","0110","0110","0111","0111"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0110","0110","0111","0110","0010","0001","0001","0001","0001","0001","0001","0100","0111","0111","0101","0011","0101","0100","0110","0100","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0011","0011","0011","0010","0011","0010","0010","0011","0011","0001","0010","0011","0010","0100","0100","0011","0001","0010","0001","0001","0010","0011","0001","0010","0010","0010","0011","0001","0010","0010","0001","0001","0010","0001","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0001","0001","0001","0001","0010","0011","0010","0010","0011","0011","0011","0010","0001","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010","0011","0011","0010","0010","0010","0001","0001","0000","0001","0001","0001","0001","0010","0010","0001","0001","0000","0000","0000","0001","0000","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0001","0001","0010","0010","0010","0011","0011","0010","0001","0110","0111","0101","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0011","0010","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0100","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0101","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0010","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0001","0001","0000","0010","0011","0011","0011","0010","0011","0100","0101","0110","0110","0010","0001","0011","1000","1000","0111","0111","1000","1000","1000","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","0111","0111","0111","0110","0101","0101","0100","0011","0011","0011","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0101","0101","0101","0100","0101","0101","0100","0100","0100","0011","0001","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0111","1000","1000","1000","1000","0111","0110","0011","0010","0010","0001","0001","0100","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0101","0111","0111","0110","0110","0111","0110"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0011","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0010","0010","0001","0001","0010","0101","0101","0110","0110","0001","0000","0000","0000","0000","0000","0000","0100","0101","0101","0101","0100","0100","0100","0101","0011","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0011","0101","0010","0100","0100","0010","0011","0100","0001","0010","0010","0010","0100","0100","0100","0010","0010","0011","0010","0001","0001","0010","0011","0010","0010","0010","0001","0011","0010","0001","0001","0010","0010","0010","0010","0011","0011","0010","0001","0001","0001","0001","0001","0010","0011","0010","0010","0010","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0001","0001","0001","0010","0001","0010","0010","0010","0001","0000","0000","0010","0011","0010","0100","0110","0110","0110","0110","0101","0101","0101","0101","0101","0010","0010","0010","0010","0010","0100","0100","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0001","0001","0001","0001","0001","0001","0001","0010","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0100","0011","0011","0100","0011","0011","0011","0011","0010","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0011","0010","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0000","0000","0000","0000","0001","0001","0001","0010","0010","0011","0010","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0101","0100","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0101","0101","0100","0101","0101","0100","0100","0101","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0010","0010","0001","0001","0001","0010","0010","0011","0011","0011","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0000","0000","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0010","0001","0011","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1000","1000","0111","0111","0101","0101","0101","0100","0010","0001","0001","0000","0001","0001","0001","0000","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0010","0100","0101","0101","0101","0101","0101","0011","0010","0110","0100","0011","0100","0001","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0011","0011","0100","0110","0111","0111","0111","0111","0101","0010","0001","0001","0001","0100","0110","0110","0110","0101","0101","0101","0101","0110","0110","0110","0110","0101","0111","0111","0110","0111","0111","0110"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0001","0010","0010","0001","0001","0010","0100","0101","0101","0101","0001","0000","0000","0000","0000","0000","0000","0100","0101","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0010","0001","0001","0001","0010","0100","0010","0011","0101","0011","0100","0011","0001","0010","0011","0011","0001","0011","0011","0010","0001","0100","0010","0001","0001","0011","0100","0010","0010","0010","0010","0100","0011","0010","0001","0001","0010","0010","0010","0010","0010","0001","0001","0011","0010","0001","0001","0010","0010","0010","0001","0001","0001","0010","0010","0010","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0000","0000","0001","0010","0011","0011","0110","1000","1000","1001","1001","1001","1001","1001","1001","1001","0110","0100","0100","0100","0101","0101","0011","0001","0010","0100","0011","0011","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0000","0001","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0001","0001","0001","0001","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0010","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0010","0011","0011","0010","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0001","0001","0010","0100","0110","0111","0111","0111","0111","0110","0110","0110","0111","0111","0111","0111","0101","0100","0010","0010","0001","0001","0001","0001","0001","0001","0000","0001","0001","0000","0000","0010","0010","0010","0010","0011","0011","0010","0001","0010","0011","0100","0011","0101","0101","0101","0101","0101","0101","0011","0011","0101","0100","0010","0100","0000","0001","0010","0010","0010","0100","0011","0100","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","0111","0111","0100","0010","0001","0001","0100","0110","0110","0101","0101","0100","0100","0101","0101","0110","0110","0101","0101","0111","0111","0110","0111","0111","0110"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0010","0010","0001","0001","0010","0100","0111","0100","0100","0001","0000","0000","0000","0000","0000","0000","0011","0100","0101","0101","0101","0011","0011","0010","0100","0101","0011","0011","0100","0010","0010","0100","0101","0011","0101","0100","0001","0011","0010","0010","0100","0010","0011","0010","0001","0010","0011","0011","0011","0100","0101","0010","0000","0011","0010","0001","0001","0011","0100","0010","0010","0001","0010","0100","0011","0010","0000","0001","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0001","0001","0000","0000","0001","0001","0010","0100","0111","1000","1000","1000","1000","1000","1000","1001","1001","0111","0100","0100","0100","0100","0101","0100","0010","0001","0011","0100","0011","0011","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0011","0010","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0001","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0000","0001","0001","0001","0010","0010","0010","0010","0001","0010","0010","0001","0010","0001","0010","0010","0010","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0010","0011","0011","0011","0100","0011","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0001","0001","0010","0010","0011","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0001","0001","0001","0001","0010","0010","0010","0001","0001","0010","0010","0001","0011","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0010","0010","0011","0010","0010","0001","0011","0010","0001","0001","0011","0011","0011","0011","0011","0010","0001","0001","0011","0101","0011","0010","0011","0011","0011","0011","0011","0010","0001","0001","0010","0010","0001","0010","0010","0010","0001","0001","0010","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0011","0011","0010","0100","0111","0101","0011","0010","0011","0101","0101","0110","0011","0001","0101","0101","0101","0101","0101","0100","0100","0100","0101","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0010","0001","0010","0010","0100","0110","0100","0011","0001","0000","0000","0000","0000","0000","0000","0011","0100","0100","0011","0100","0011","0100","0011","0110","0110","0101","0011","0010","0010","0010","0100","0101","0100","0101","0101","0010","0011","0011","0011","0100","0010","0010","0010","0001","0010","0011","0011","0101","0101","0110","0101","0010","0010","0010","0000","0010","0100","0100","0001","0001","0001","0001","0010","0001","0000","0000","0000","0001","0010","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0000","0000","0001","0001","0001","0010","0100","0110","0111","0111","0111","0111","0111","1000","1000","1000","0101","0011","0100","0100","0100","0101","0100","0001","0001","0011","0100","0011","0011","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0100","0011","0100","0100","0011","0100","0100","0011","0011","0001","0000","0000","0000","0000","0000","0001","0010","0011","0011","0011","0100","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0001","0010","0010","0011","0010","0010","0001","0010","0010","0001","0001","0001","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0010","0010","0010","0011","0011","0010","0100","0011","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0011","0010","0010","0001","0001","0001","0010","0010","0011","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0001","0010","0010","0100","0101","0101","0101","0011","0010","0010","0001","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0100","0100","0011","0011","0100","0100","0100","0101","0110","0101","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0011","0011","0010","0011","0101","0110","0100","0011","0011","0011","0100","0100","0101","0101","0101","0101","0101","0101","0100","0011","0100","0101","0101","0101","0101","0101","0110","0110","0111","0111","0111","0101"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0100","0011","0011","0011","0010","0011","0011","0011","0011","0010","0101","0111","0101","0011","0001","0000","0000","0000","0000","0000","0000","0010","0101","0011","0011","0011","0011","0100","0011","0101","0111","0101","0101","0100","0100","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0001","0001","0001","0001","0010","0011","0011","0100","0100","0100","0100","0011","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0000","0001","0001","0001","0010","0010","0010","0010","0011","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0000","0000","0000","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0101","0101","0011","0001","0001","0011","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0010","0010","0001","0001","0001","0001","0001","0010","0010","0011","0011","0011","0010","0010","0011","0010","0011","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0000","0000","0001","0001","0010","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0011","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0011","0010","0010","0100","0010","0010","0011","0100","0100","0011","0010","0010","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0010","0010","0010","0011","0010","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0001","0001","0001","0001","0001","0010","0011","0101","0101","0101","0101","0100","0011","0011","0101","0101","0110","0110","0110","0101","0110","0111","0111","0111","0110"),
("0100","0010","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0111","0111","0101","0011","0011","0100","0100","0101","0111","0111","0111","0111","0110","0111","0110","0110","0110","0110","0111","0110","0101","0110","0100","0011","0011","0011","0100","0100","0011","0101","0110","0101","0101","0010","0000","0000","0000","0000","0000","0000","0010","0100","0011","0100","0101","0011","0100","0011","0010","0101","0101","0100","0011","0100","0101","0011","0001","0010","0011","0010","0011","0100","0011","0110","0101","0001","0010","0010","0001","0001","0001","0000","0000","0000","0001","0000","0000","0000","0010","0010","0001","0001","0010","0010","0001","0001","0001","0000","0000","0000","0001","0001","0000","0000","0000","0001","0001","0010","0011","0010","0001","0010","0001","0001","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0000","0000","0000","0000","0000","0001","0000","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0010","0000","0010","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0100","0011","0011","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0101","0100","0011","0011","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0011","0011","0100","0010","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0100","0011","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0011","0011","0010","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0001","0001","0001","0001","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0011","0010","0001","0000","0001","0001","0001","0001","0010","0001","0101","0110","0011","0010","0001","0001","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0010","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0001","0010","0010","0010","0011","0010","0011","0011","0010","0011","0010","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0010","0011","0011","0100","0100","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0101","0100","0011","0100","0011","0010","0001","0001","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0101","0101","0101","0101","0011","0011","0011","0101","0101","0101","0110","0110","0101","0111","0111","0111","0111","0101"),
("0110","0011","1000","1001","0111","0011","0111","1000","0111","0010","0110","0111","0110","0010","0101","0111","0110","0011","0101","0111","1000","0101","0000","0000","0000","0000","0011","1000","0111","0111","1000","0111","0100","0001","0001","0001","0011","0111","0111","0110","0110","0110","0100","0011","0010","0010","0010","0010","0101","0101","0011","0101","0001","0000","0000","0000","0000","0000","0000","0011","0100","0100","0100","0100","0100","0100","0010","0001","0011","0101","0100","0011","0010","0101","0101","0011","0010","0101","0100","0100","0011","0010","0100","0100","0010","0001","0010","0001","0001","0001","0000","0000","0000","0001","0000","0000","0000","0011","0011","0001","0011","0011","0010","0001","0010","0001","0000","0001","0001","0000","0001","0000","0000","0001","0011","0011","0011","0011","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0001","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0000","0000","0001","0000","0000","0000","0000","0010","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0100","0011","0011","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0101","0100","0100","0100","0011","0010","0011","0010","0010","0011","0011","0010","0010","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0010","0010","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0010","0011","0100","0011","0100","0100","0011","0011","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0010","0001","0010","0010","0001","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0101","0100","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0010","0010","0011","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0001","0001","0001","0001","0011","0101","0100","0110","0101","0001","0001","0001","0001","0010","0100","0101","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0100","0101","0101","0011","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0000","0000","0001","0000","0001","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0101","0110","0110","0101","0011","0010","0011","0101","0101","0101","0110","0110","0101","0110","0110","0111","0111","0101"),
("0010","0111","1010","1001","0100","0110","1001","1001","0100","0110","1001","1001","0100","0101","1001","1001","0101","0010","0110","1000","1000","0101","0001","0001","0010","0010","0100","1000","1000","1000","0111","1000","0101","0001","0001","0001","0011","0110","0111","0111","0101","0110","0110","0010","0000","0000","0000","0000","0011","0100","0011","0101","0010","0000","0000","0000","0000","0000","0000","0100","0100","0100","0011","0011","0011","0100","0011","0010","0010","0011","0100","0010","0010","0011","0011","0101","0010","0011","0011","0101","0100","0001","0011","0101","0001","0010","0011","0001","0010","0011","0000","0000","0000","0000","0000","0000","0000","0100","0011","0001","0011","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0011","0010","0010","0100","0011","0001","0010","0010","0001","0001","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0000","0001","0000","0001","0001","0001","0001","0010","0010","0010","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0101","0100","0100","0101","0100","0011","0100","0011","0010","0010","0010","0011","0010","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0100","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0011","0011","0100","0100","0011","0100","0011","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0010","0001","0001","0010","0010","0010","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0010","0001","0001","0010","0010","0011","0101","0101","0110","0101","0001","0001","0000","0001","0001","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0100","0100","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0101","0110","0110","0101","0100","0011","0011","0101","0101","0110","0110","0110","0101","0110","0111","0111","0110","0101"),
("0110","1010","1010","0101","0101","1001","1001","0101","0100","1001","1001","0101","0011","1000","1001","0101","0010","0011","0110","1000","1000","0110","0001","0001","0010","0010","0100","1000","1000","1000","1000","0111","0110","0001","0001","0010","0100","0111","1000","0111","0110","0101","0110","0010","0000","0001","0001","0001","0011","0100","0101","0101","0010","0000","0000","0000","0000","0000","0000","0010","0011","0010","0100","0011","0100","0100","0011","0001","0010","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0100","0101","0010","0101","0100","0001","0100","0100","0001","0011","0100","0000","0000","0000","0000","0000","0000","0000","0010","0010","0001","0010","0010","0010","0010","0001","0010","0001","0000","0001","0000","0001","0010","0011","0010","0010","0011","0010","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0001","0001","0001","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0011","0010","0001","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0001","0000","0001","0001","0001","0011","0100","0100","0011","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0010","0001","0001","0010","0001","0001","0010","0001","0010","0011","0011","0011","0100","0011","0011","0100","0100","0011","0100","0011","0011","0100","0011","0100","0101","0100","0100","0101","0100","0100","0101","0100","0100","0101","0100","0100","0101","0011","0010","0010","0001","0010","0011","0011","0100","0101","0100","0100","0100","0011","0100","0100","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0010","0010","0010","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0011","0011","0100","0101","0010","0010","0010","0010","0001","0010","0101","0101","0110","0101","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0100","0110","0011","0000","0010","0010","0001","0001","0001","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0001","0001","0001","0001","0001","0001","0011","0001","0000","0001","0001","0001","0001","0001","0001","0001","0011","0101","0110","0101","0101","0101","0101","0101","0101","0110","0110","0110","0111","0110","0111","0111","0111","0111","0101"),
("1001","1010","0110","0100","1001","1010","0110","0011","1000","1001","0110","0011","0111","1001","0111","0010","0010","0011","0110","1000","1000","0110","0001","0001","0011","0011","0101","1000","1000","1000","0111","0110","0110","0001","0001","0010","0100","1000","1000","1000","0111","0101","0100","0011","0000","0001","0001","0001","0010","0011","0110","0101","0010","0000","0000","0000","0000","0000","0000","0010","0100","0101","0011","0100","0011","0100","0100","0010","0000","0000","0000","0000","0000","0001","0001","0000","0000","0001","0010","0010","0110","0100","0001","0001","0010","0100","0101","0010","0010","0011","0001","0001","0000","0000","0000","0000","0000","0100","0011","0000","0001","0010","0001","0010","0010","0010","0001","0000","0000","0000","0000","0000","0000","0001","0011","0011","0010","0001","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0011","0100","0100","0011","0011","0011","0011","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0010","0011","0100","0011","0011","0011","0011","0011","0010","0010","0001","0001","0001","0001","0010","0001","0001","0000","0000","0000","0001","0011","0011","0011","0100","0100","0011","0100","0100","0011","0011","0011","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0100","0011","0011","0100","0100","0011","0100","0100","0011","0100","0100","0100","0101","0100","0100","0101","0100","0100","0101","0100","0100","0101","0100","0100","0101","0100","0100","0100","0010","0010","0011","0010","0011","0101","0100","0100","0101","0100","0100","0101","0100","0011","0100","0100","0011","0100","0100","0011","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0011","0011","0011","0010","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0010","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0100","0101","0101","0111","0011","0010","0010","0001","0000","0001","0100","0101","0110","0101","0001","0010","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0011","0100","0011","0011","0001","0000","0000","0000","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0001","0011","0001","0000","0000","0001","0001","0001","0001","0001","0000","0011","0101","0110","0110","0110","0110","0101","0110","0101","0110","0110","0110","0111","0110","0111","0111","0111","0110","0101"),
("0111","0110","0010","0110","0111","0110","0011","0110","1000","0111","0011","0110","1000","0111","0010","0010","0010","0011","0110","1001","1000","0110","0001","0001","0011","0011","0101","1000","1001","1001","1000","0111","0110","0010","0001","0001","0011","0111","0111","1000","0111","0110","0100","0010","0000","0001","0001","0001","0010","0011","0100","0101","0010","0000","0000","0000","0000","0000","0000","0011","0100","0100","0010","0010","0010","0100","0101","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","0011","0110","0011","0000","0010","0010","0011","0110","0010","0010","0010","0001","0000","0000","0000","0000","0000","0000","0010","0010","0001","0001","0010","0001","0001","0001","0010","0001","0000","0000","0000","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0100","0100","0100","0100","0011","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0010","0001","0010","0010","0010","0011","0011","0011","0010","0010","0001","0000","0000","0000","0001","0010","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0010","0011","0010","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0100","0011","0101","0100","0011","0101","0100","0011","0101","0100","0100","0101","0100","0100","0101","0100","0100","0101","0100","0100","0101","0011","0011","0011","0011","0011","0100","0100","0100","0101","0100","0100","0101","0100","0011","0100","0100","0011","0100","0011","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0001","0010","0011","0011","0011","0011","0010","0010","0001","0001","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0011","0010","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0100","0101","0101","0110","0010","0001","0001","0001","0000","0001","0100","0101","0110","0101","0100","0110","0111","0111","0011","0010","0010","0010","0011","0010","0011","0010","0011","0010","0011","0011","0011","0011","0011","0010","0010","0010","0011","0100","0001","0000","0000","0000","0000","0000","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0001","0000","0000","0001","0001","0001","0001","0001","0000","0011","0101","0101","0110","0101","0110","0101","0100","0011","0011","0011","0101","0111","0110","0111","0111","0111","0110","0101"),
("0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0010","0010","0010","0011","0011","0101","1000","1001","0111","0010","0010","0011","0011","0100","1000","1001","1001","1000","0111","0110","0010","0010","0010","0010","0111","0111","1000","0111","0111","0101","0011","0000","0001","0001","0001","0010","0011","0101","0110","0010","0000","0000","0000","0000","0000","0000","0001","0011","0100","0010","0011","0010","0010","0011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0010","0101","0010","0000","0010","0010","0011","0011","0001","0010","0010","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0000","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0100","0011","0011","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0100","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0010","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0011","0100","0100","0011","0011","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0010","0001","0010","0010","0001","0010","0001","0001","0001","0001","0001","0011","0011","0100","0100","0010","0010","0011","0011","0011","0011","0011","0010","0010","0001","0000","0000","0000","0000","0000","0000","0010","0011","0010","0001","0010","0010","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0011","0100","0011","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0101","0100","0100","0101","0100","0011","0100","0011","0011","0100","0011","0011","0100","0100","0011","0101","0100","0011","0100","0100","0011","0100","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0010","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0011","0010","0001","0001","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0100","0101","0110","0110","0010","0000","0000","0000","0000","0000","0011","0100","0110","0110","0111","0111","0111","0111","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0011","0011","0010","0001","0001","0001","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0010","0001","0010","0001","0001","0001","0001","0010","0010","0011","0101","0101","0110","0110","0110","0101","0000","0000","0000","0001","0101","0110","0110","0111","0111","0110","0110","0100"),
("0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0100","0011","0111","0111","0111","0010","0010","0011","0011","0100","1000","1000","1000","1000","0111","0101","0001","0010","0011","0011","0101","0101","0111","0111","0110","0111","0100","0000","0001","0001","0001","0001","0010","0101","0110","0010","0001","0001","0000","0000","0000","0000","0001","0100","0101","0011","0011","0010","0001","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0011","0011","0001","0011","0010","0001","0010","0011","0001","0010","0010","0000","0001","0000","0000","0001","0000","0000","0000","0000","0001","0010","0010","0011","0010","0000","0001","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0011","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0100","0011","0011","0011","0101","0011","0001","0000","0001","0001","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0100","0011","0010","0100","0100","0011","0011","0010","0010","0001","0000","0000","0000","0001","0001","0001","0010","0011","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0011","0010","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0010","0001","0001","0001","0000","0000","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0001","0001","0100","0101","0101","0111","0010","0001","0001","0001","0011","0011","0011","0100","0110","0111","0111","0111","0111","0111","0101","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","0100","0100","0011","0001","0001","0001","0001","0001","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0100","0100","0011","0011","0011","0100","0011","0100","0100","0011","0011","0100","0011","0100","0100","0100","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0110","0110","0110","0110","0110","0101","0000","0000","0000","0001","0101","0110","0110","0110","0110","0110","0101","0100"),
("0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0011","0011","0110","0110","0110","0100","0100","0011","0011","0100","1000","1000","0111","0111","0110","0101","0001","0001","0010","0011","0110","0101","0100","0110","0101","0101","0101","0001","0001","0001","0001","0010","0010","0110","0101","0101","0110","0101","0001","0001","0001","0000","0001","0011","0011","0011","0011","0100","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0011","0010","0001","0011","0010","0001","0010","0010","0001","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0010","0001","0010","0010","0011","0001","0001","0000","0000","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0000","0000","0001","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0011","0011","0010","0010","0010","0001","0001","0001","0001","0001","0011","0011","0010","0011","0011","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0100","0011","0011","0100","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0100","0011","0011","0010","0011","0011","0011","0100","0011","0011","0011","0011","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0010","0001","0011","0011","0010","0011","0100","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0010","0010","0011","0100","0101","0011","0000","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0011","0010","0010","0001","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0001","0000","0000","0000","0000","0000","0001","0001","0010","0010","0010","0010","0011","0011","0011","0010","0011","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0001","0001","0100","0101","0101","0111","0011","0010","0100","0101","0110","0101","0011","0100","0101","0110","0111","1000","0111","0111","0101","0100","0011","0100","0100","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0001","0001","0000","0001","0001","0010","0011","0011","0011","0011","0011","0011","0010","0000","0001","0010","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0101","0101","0101","0101","0110","0110","0101","0011","0010","0010","0010","0011","0100","0011","0100","0100","0100","0011","0100","0101","0110","0110","0110","0110","0101","0001","0000","0001","0010","0101","0110","0110","0110","0110","0110","0110","0101"),
("0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0110","0011","0010","0011","0010","0011","0100","0100","0110","0110","0110","0111","0111","0111","0110","0111","0110","0101","0010","0001","0001","0011","0101","0101","0100","0100","0100","0011","0011","0010","0010","0001","0010","0010","0010","0100","0110","0111","0110","0101","0001","0000","0001","0001","0010","0010","0010","0001","0001","0010","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0100","0001","0001","0011","0010","0001","0011","0011","0001","0010","0011","0001","0000","0000","0000","0000","0000","0000","0000","0011","0011","0001","0001","0010","0100","0010","0000","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0000","0000","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0011","0011","0010","0011","0011","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0011","0100","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0011","0010","0001","0011","0010","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0011","0100","0100","0101","0101","0101","0011","0000","0000","0001","0010","0010","0011","0011","0011","0100","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0010","0010","0010","0010","0011","0100","0011","0100","0101","0010","0001","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0000","0000","0011","0101","0101","0111","0110","0110","0111","0111","0111","0101","0011","0100","0100","0110","0111","0111","0111","0111","0101","0100","0100","0110","0110","0110","0110","0110","0110","0110","0101","0011","0100","0100","0101","0100","0011","0011","0100","0101","0100","0010","0001","0001","0001","0001","0001","0010","0010","0011","0011","0011","0011","0010","0001","0001","0010","0011","0011","0011","0011","0011","0010","0001","0001","0001","0010","0010","0001","0001","0001","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0001","0010","0010","0011","0100","0011","0010","0011","0011","0011","0011","0011","0011","0010","0000","0000","0001","0010","0100","0101","0100","0101","0101","0110","0101","0011"),
("0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0110","0100","0001","0001","0010","0001","0010","0100","0100","0101","0110","0110","0111","0111","0111","0101","0110","0111","0100","0001","0001","0001","0011","0111","0101","0101","0100","0001","0010","0010","0010","0100","0001","0010","0011","0010","0011","0100","0110","0110","0100","0001","0000","0000","0000","0010","0011","0011","0011","0010","0001","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0011","0011","0001","0010","0011","0010","0011","0001","0000","0011","0100","0001","0000","0000","0000","0000","0000","0000","0001","0011","0011","0001","0001","0010","0011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0000","0000","0001","0001","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0100","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0101","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0101","0101","0101","0101","0101","0011","0010","0001","0001","0010","0010","0011","0010","0010","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0100","0101","0101","0101","0101","0101","0101","0110","0101","0001","0000","0001","0001","0010","0011","0011","0010","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0001","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0000","0001","0001","0000","0000","0000","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0100","0100","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0000","0000","0000","0001","0011","0100","0100","0111","0111","0111","0111","0111","0111","0101","0100","0100","0100","0111","0111","0111","0111","0111","0110","0101","0100","0101","0110","0101","0110","0101","0110","0100","0011","0101","0110","0101","0101","0100","0010","0011","0110","0110","0101","0010","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0000","0000","0000","0001","0001","0010","0011","0011","0011","0010","0011","0100","0011"),
("0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0100","0100","0001","0000","0001","0001","0001","0010","0011","0010","0011","0100","0101","0101","0101","0101","0101","0100","0110","0101","0001","0001","0010","0010","0101","0100","0011","0010","0001","0001","0001","0001","0010","0001","0000","0001","0001","0010","0011","0101","0100","0100","0000","0000","0000","0000","0010","0100","0011","0011","0011","0010","0001","0010","0001","0000","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","0011","0011","0001","0010","0010","0001","0011","0001","0001","0010","0010","0001","0000","0001","0001","0001","0000","0000","0000","0010","0011","0010","0001","0010","0010","0010","0010","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0010","0001","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0001","0001","0001","0010","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0100","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0100","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0101","0011","0010","0001","0001","0001","0011","0100","0011","0010","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0010","0000","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0010","0010","0011","0011","0011","0110","0110","0011","0010","0010","0010","0001","0001","0001","0000","0000","0001","0001","0010","0100","0100","0011","0100","0100","0111","0111","0111","0111","0111","0111","0101","0011","0011","0100","0110","0111","0111","0111","0111","0110","0101","0100","0101","0101","0101","0110","0101","0101","0011","0010","0011","0101","0110","0110","0111","0110","0101","0100","0011","0011","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0001","0001","0011","0100","0101","0100","0011","0011","0100","0100"),
("0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0100","0100","0101","0101","0101","0100","0101","0101","0001","0001","0001","0010","0101","0101","0011","0010","0001","0001","0001","0001","0001","0000","0000","0001","0010","0010","0011","0101","0100","0011","0001","0000","0000","0000","0010","0101","0010","0011","0011","0001","0000","0001","0001","0000","0000","0001","0010","0001","0000","0001","0001","0001","0001","0010","0011","0011","0001","0001","0010","0001","0010","0010","0010","0011","0010","0001","0001","0001","0001","0001","0001","0000","0000","0010","0011","0010","0001","0001","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0001","0000","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0000","0000","0000","0000","0000","0001","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0111","1000","1000","1000","1000","1000","1000","1000","0111","0111","1000","0111","0111","0111","0111","0111","0110","0101","0011","0010","0010","0011","0100","0100","0011","0010","0001","0001","0000","0001","0011","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0000","0001","0001","0001","0010","0011","0010","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0010","0011","0100","0011","0011","0100","0010","0011","0011","0010","0011","0011","0011","0011","0100","0010","0011","0011","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0010","0001","0001","0001","0010","0100","0100","0100","0111","0110","0010","0010","0001","0001","0001","0000","0000","0001","0010","0011","0101","0110","0110","0101","0011","0100","0100","0111","0111","0111","0111","1000","0111","0101","0011","0011","0011","0101","0111","0111","0111","0111","0110","0101","0100","0101","0101","0110","0101","0101","0011","0010","0011","0100","0101","0110","0110","0110","0100","0100","0011","0011","0011","0010","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011"),
("0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0010","0001","0001","0001","0001","0000","0000","0001","0001","0001","0010","0100","0011","0010","0001","0000","0000","0000","0001","0011","0010","0010","0011","0011","0010","0010","0011","0010","0000","0001","0010","0001","0000","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0000","0001","0001","0010","0010","0001","0000","0001","0011","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0001","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0011","0010","0011","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0110","0101","0100","0010","0010","0011","0101","0110","0110","0101","0110","0110","0110","0101","0011","0010","0001","0001","0001","0011","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","1000","0111","0111","1000","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0100","0000","0000","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0001","0001","0000","0000","0000","0000","0000","0001","0000","0001","0001","0001","0001","0010","0010","0100","0100","0100","0101","0110","0001","0001","0000","0000","0001","0001","0010","0100","0101","0110","0111","0111","0111","0110","0011","0100","0011","0110","0111","0111","0111","0110","0101","0111","0110","0011","0100","0110","0111","0111","0111","0111","0101","0100","0100","0101","0101","0101","0101","0100","0010","0010","0011","0011","0101","0110","0111","0100","0010","0100","0110","0101","0101","0001","0001","0001","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0100","0011","0011","0011","0100","0100","0001","0000","0001","0010","0010","0010","0001","0001","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010"),
("0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0011","0010","0001","0011","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0010","0010","0010","0011","0100","0100","0011","0011","0100","0011","0001","0000","0001","0001","0001","0001","0010","0010","0010","0001","0000","0000","0000","0001","0010","0010","0100","0100","0101","0101","0011","0011","0110","0010","0000","0000","0001","0000","0001","0001","0010","0010","0001","0001","0001","0001","0000","0001","0001","0010","0001","0001","0011","0011","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0011","0101","0101","0101","0101","0101","0101","0100","0101","0010","0001","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0000","0001","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0010","0011","0011","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0101","0100","0010","0010","0011","0101","0110","0110","0101","0111","0100","0011","0100","0011","0100","0111","0110","0110","0100","0010","0001","0001","0001","0010","0011","0101","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0110","0110","0110","0101","0001","0000","0001","0001","0010","0010","0010","0010","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0010","0001","0010","0001","0010","0100","0100","0100","0100","0110","0001","0000","0001","0010","0011","0100","0101","0110","0111","0110","0111","0111","0111","0110","0011","0100","0011","0110","0111","0111","0111","0100","0100","0111","0101","0011","0100","0110","0111","0111","0111","0111","0101","0100","0011","0100","0101","0101","0011","0001","0001","0001","0011","0100","0100","0101","0101","0100","0101","0101","0101","0101","0110","0101","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0100","0010","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0011","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010"),
("0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0100","0111","0111","0111","0110","0110","0110","0110","0110","0110","0111","0111","0110","0101","0101","0111","0110","0110","0101","0100","0010","0010","0001","0001","0010","0100","0101","0011","0011","0011","0011","0011","0010","0011","0001","0000","0010","0001","0001","0010","0011","0001","0000","0000","0000","0001","0011","0010","0011","0011","0011","0101","0101","0010","0011","0010","0010","0000","0000","0000","0001","0010","0010","0011","0001","0001","0001","0010","0001","0000","0001","0001","0001","0001","0010","0001","0000","0000","0000","0000","0001","0001","0001","0001","0000","0001","0001","0000","0000","0000","0011","0101","0101","0101","0101","0101","0101","0101","0101","0011","0001","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0010","0000","0000","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0010","0100","0011","0010","0011","0011","0011","0011","0011","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1000","1000","1000","1000","1000","0111","0111","0110","0100","0011","0010","0010","0011","0101","0110","0110","0101","0110","0100","0011","0101","0100","0100","0100","0011","0100","0110","0100","0101","0111","0110","0101","0100","0010","0001","0000","0001","0010","0100","0110","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0110","0010","0100","0110","0001","0000","0001","0001","0001","0010","0010","0010","0011","0011","0010","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0010","0001","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0011","0100","0100","0100","0101","0001","0010","0011","0101","0110","0110","0111","0111","0111","0111","0111","0110","0110","0110","0011","0011","0011","0110","0111","0111","0111","0011","0011","0111","0101","0011","0100","0110","0111","0111","0111","0111","0110","0101","0100","0101","0101","0100","0010","0001","0010","0001","0001","0010","0011","0011","0001","0010","0011","0101","0110","1000","1000","1000","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0010","0001","0001","0010","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0001"),
("0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0011","0010","0011","0111","0111","0110","0011","0001","0001","0010","0010","0101","0111","0111","0111","0111","0101","0100","0100","0011","0100","0100","0010","0100","0001","0001","0011","0100","0100","0101","0100","0011","0010","0011","0010","0011","0010","0001","0001","0001","0010","0010","0011","0001","0000","0000","0000","0001","0101","0101","0011","0010","0001","0011","0011","0010","0001","0010","0011","0011","0001","0001","0001","0001","0010","0011","0010","0010","0001","0010","0010","0000","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0001","0001","0000","0100","0101","0101","0110","0110","0101","0101","0101","0101","0011","0001","0100","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0111","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0011","0000","0000","0001","0010","0010","0010","0011","0011","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0100","0011","0010","0011","0011","0010","0011","0011","0011","0110","0110","0110","0110","0111","0111","0111","0110","0111","0110","0101","1000","1000","0111","0111","0110","0100","0011","0010","0010","0100","0101","0110","0110","0101","0110","0100","0011","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0101","0101","0111","0110","0101","0011","0001","0000","0000","0001","0011","0101","0111","0111","1000","1000","1000","1000","1000","1000","0111","0110","0110","0110","0111","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0010","0011","0011","0000","0001","0001","0001","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0100","0011","0100","0100","0011","0011","0100","0011","0011","0100","0011","0100","0100","0011","0011","0011","0011","0011","0100","0010","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0011","0100","0011","0100","0110","0100","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110","0101","0110","0101","0011","0011","0010","0101","0110","0111","0111","0011","0010","0110","0101","0011","0100","0110","0111","0111","0111","0111","0110","0101","0100","0101","0101","0011","0010","0011","0011","0011","0011","0100","0100","0010","0010","0101","0110","0101","0101","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0001","0010","0010","0010"),
("0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0001","0010","0010","0011","0111","0111","0111","0011","0000","0000","0000","0000","0101","0111","0101","0110","1000","0111","0010","0000","0000","0000","0000","0010","0100","0001","0010","0011","0011","0001","0001","0001","0001","0001","0001","0011","0010","0010","0001","0001","0011","0011","0101","0011","0000","0000","0000","0000","0011","0101","0011","0010","0010","0100","0100","0100","0010","0010","0010","0010","0011","0010","0001","0001","0001","0010","0001","0010","0010","0011","0100","0101","0010","0000","0010","0001","0001","0001","0001","0001","0000","0000","0000","0001","0000","0001","0001","0001","0001","0000","0000","0001","0001","0011","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0001","0101","0110","0101","0010","0100","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0100","0011","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0110","0111","0110","0111","0111","0111","0111","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0100","0011","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0100","0101","0101","0100","0011","0010","0011","0100","0110","0110","0110","0101","0110","0100","0011","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0100","0100","0110","0110","0101","0110","0110","0100","0010","0001","0000","0001","0010","0011","0101","0111","1000","1000","1000","1000","0111","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0011","0001","0000","0000","0001","0001","0010","0010","0010","0010","0011","0010","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0010","0010","0010","0010","0011","0001","0001","0001","0001","0001","0010","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0000","0010","0100","0011","0100","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0101","0011","0011","0011","0101","0110","0111","0111","0011","0011","0100","0011","0011","0011","0101","0111","0111","0111","0111","0110","0101","0100","0101","0100","0011","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0101","0100","0001","0010","0001","0001","0001","0001","0001"),
("0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0001","0010","0010","0011","0111","0111","0111","0011","0000","0000","0000","0000","0101","0111","0101","0111","1000","0111","0100","0000","0000","0000","0000","0010","0101","0001","0011","0100","0011","0001","0000","0000","0000","0000","0010","0100","0011","0011","0011","0001","0110","0110","0011","0010","0000","0000","0000","0001","0010","0100","0100","0011","0001","0010","0101","0010","0010","0011","0010","0001","0010","0100","0001","0001","0001","0001","0011","0010","0010","0001","0010","0100","0010","0001","0100","0001","0000","0010","0010","0001","0000","0001","0001","0001","0000","0001","0001","0000","0001","0010","0011","0011","0100","0011","0001","0001","0001","0001","0001","0001","0010","0001","0001","0000","0000","0001","0010","0010","0000","0001","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0111","0100","0010","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0000","0000","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0011","0010","0011","0011","0010","0011","0011","0110","0110","0110","0110","0110","0110","0110","0110","0100","0011","0001","0001","0001","0011","0100","0110","0110","0110","0101","0110","0100","0011","0101","0100","0100","0100","0100","0100","0101","0101","0011","0011","0100","0100","0100","0100","0100","0101","0101","0100","0100","0100","0101","0101","0101","0100","0110","0110","0101","0110","0101","0011","0001","0001","0000","0001","0010","0100","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0111","0101","0001","0000","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0010","0011","0011","0100","0110","0110","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0101","0011","0100","0011","0110","0111","0111","0111","0100","0101","0100","0010","0010","0100","0110","0111","0111","0111","0111","0110","0100","0100","0100","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","0101","0101","0110","0101","0001","0010","0001","0001","0001","0001","0001"),
("0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0010","0010","0011","0111","0111","0111","0100","0000","0000","0000","0000","0101","0111","0110","0110","0111","0110","0100","0001","0000","0000","0000","0010","0011","0001","0100","0100","0100","0100","0001","0000","0000","0000","0000","0001","0010","0011","0011","0001","0100","0111","0101","0010","0000","0000","0000","0000","0001","0011","0011","0100","0010","0010","0100","0011","0010","0000","0000","0000","0001","0001","0001","0001","0001","0000","0000","0010","0101","0011","0010","0010","0010","0010","0011","0001","0001","0011","0011","0001","0000","0001","0001","0001","0000","0001","0010","0000","0001","0010","0011","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0111","0111","0111","0110","0010","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0010","0000","0000","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0110","0110","0110","0110","0110","0101","0100","0010","0001","0001","0011","0011","0011","0110","0110","0101","0110","0100","0011","0100","0100","0100","0100","0100","0100","0101","0101","0110","0110","0110","0010","0001","0000","0000","0000","0000","0001","0001","0000","0001","0000","0011","0110","0110","0101","0101","0101","0101","0100","0110","0111","0110","0101","0100","0011","0001","0001","0001","0001","0011","0100","0110","1000","1000","1001","1001","1001","1001","1001","1001","1001","1000","0111","0110","0110","0110","0010","0000","0001","0001","0001","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0100","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0100","0011","0011","0011","0010","0001","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0000","0000","0000","0010","0011","0011","0100","0110","0110","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0110","0110","0101","0011","0011","0011","0110","0111","0111","0111","0101","0110","0100","0011","0011","0100","0110","0111","0111","0111","0111","0101","0100","0010","0011","0010","0001","0001","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0100","0101","0101","0110","0110","0100","0001","0001","0010","0010","0001","0001","0001"),
("0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0011","0010","0011","0111","0111","0111","0100","0000","0000","0000","0000","0101","0111","0110","0101","0110","0110","0100","0001","0000","0000","0000","0001","0011","0010","0100","0101","0110","0100","0001","0000","0000","0000","0001","0010","0010","0010","0100","0010","0011","0100","0100","0011","0001","0000","0001","0000","0001","0011","0010","0100","0010","0001","0010","0011","0010","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0100","0110","0011","0011","0001","0001","0010","0010","0001","0010","0010","0001","0000","0001","0001","0001","0001","0001","0001","0001","0010","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0000","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0011","0110","0110","0110","0101","0100","0010","0010","0010","0100","0101","0110","0101","0011","0101","0011","0011","0100","0100","0100","0100","0100","0100","0101","0101","0110","0110","0110","0110","0111","0110","0011","0010","0000","0000","0000","0000","0010","0011","0000","0001","0001","0011","0111","0110","0110","0110","0101","0101","0101","0101","0101","0100","0110","0111","0110","0100","0010","0001","0001","0000","0001","0001","0010","0100","0110","0110","0110","0110","0110","0111","0111","0110","0110","0110","0110","0011","0000","0001","0001","0001","0010","0010","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0100","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0000","0001","0001","0001","0010","0011","0010","0010","0011","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0000","0000","0000","0001","0010","0010","0010","0011","0100","0100","0000","0000","0001","0010","0011","0011","0100","0110","0110","0111","0111","0111","0111","0111","0111","0101","0101","1000","0111","0111","0111","0101","0011","0100","0011","0110","0111","0111","0111","0110","0110","0100","0011","0011","0100","0111","0111","0111","0111","0111","0101","0011","0011","0101","0100","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0000","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0001","0100","0100","0011","0101","0110","0100","0001","0001","0010","0010","0010","0010","0001"),
("0100","0011","0101","0101","0101","0100","0101","0101","0110","0101","0101","0101","0011","0011","0011","0111","0111","0111","0100","0000","0000","0000","0000","0101","0111","0110","0110","0110","0101","0011","0000","0001","0000","0000","0010","0101","0010","0100","0110","0110","0100","0001","0000","0000","0000","0001","0100","0100","0100","0011","0001","0011","0101","0101","0011","0001","0000","0000","0000","0001","0101","0011","0100","0101","0010","0010","0011","0010","0000","0001","0001","0000","0001","0001","0000","0001","0001","0001","0001","0010","0100","0011","0010","0001","0000","0010","0010","0001","0001","0011","0001","0000","0000","0000","0000","0001","0001","0010","0001","0010","0011","0010","0100","0011","0100","0100","0011","0101","0011","0100","0100","0011","0101","0100","0011","0010","0100","0011","0100","0101","0011","0101","0100","0100","0101","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0010","0100","0100","0011","0010","0011","0100","0101","0110","0101","0110","0100","0011","0011","0100","0100","0100","0100","0100","0100","0101","0101","0110","0110","0110","0110","0111","0111","0111","0111","0111","0011","0010","0001","0000","0000","0000","0010","0011","0000","0001","0010","0011","0111","0111","0111","0111","0110","0110","0110","0101","0101","0100","0101","0101","0100","0101","0101","0100","0011","0001","0000","0000","0000","0010","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0100","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0010","0011","0011","0010","0011","0011","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0011","0100","0011","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0011","0011","0010","0010","0010","0011","0011","0011","0011","0010","0010","0001","0001","0000","0000","0000","0000","0001","0010","0010","0011","0100","0101","0101","0110","0101","0000","0000","0001","0011","0011","0011","0100","0101","0110","0111","0111","0111","0111","0111","0111","0100","0100","0110","0101","0111","0111","0101","0100","0100","0011","0101","0110","0111","0111","0111","0110","0100","0011","0011","0101","0111","0111","0111","0111","0111","0101","0100","0101","0101","0101","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0001","0001","0010","0010","0001","0010","0010","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0100","0100","0011","0100","0101","0010","0001","0001","0001","0010","0010","0010","0010"),
("0011","0100","0011","0011","0010","0011","0010","0100","0101","0110","0101","0101","0100","0011","0011","0110","0111","0111","0100","0000","0000","0000","0000","0101","0111","0111","0111","0110","0110","0011","0001","0001","0000","0000","0010","0100","0011","0101","0110","0111","0100","0001","0000","0000","0000","0001","0010","0011","0100","0011","0010","0001","0101","0100","0010","0001","0000","0000","0010","0001","0100","0100","0101","0101","0011","0010","0010","0010","0000","0001","0010","0001","0001","0010","0001","0000","0000","0000","0001","0001","0011","0010","0010","0010","0000","0011","0011","0001","0010","0011","0001","0000","0000","0000","0000","0001","0001","0001","0001","0010","0011","0001","0001","0010","0011","0011","0011","0100","0011","0100","0100","0011","0100","0010","0001","0011","0100","0011","0100","0100","0011","0100","0100","0011","0101","0011","0011","0101","0010","0100","0100","0010","0100","0100","0011","0101","0011","0011","0101","0011","0100","0100","0011","0101","0100","0011","0101","0100","0100","0101","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0011","0100","0101","0110","0110","0110","0100","0010","0100","0011","0011","0011","0100","0100","0100","0101","0101","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0011","0010","0001","0000","0000","0000","0010","0011","0000","0001","0001","0011","0111","0111","0111","0111","0111","0111","0110","0110","0110","0101","0101","0100","0100","0101","0110","0101","0110","0101","0011","0010","0001","0000","0001","0010","0100","0101","0110","0110","0110","0110","0110","0101","0001","0000","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0010","0011","0100","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0001","0001","0001","0000","0001","0001","0001","0010","0010","0010","0011","0100","0101","0110","0110","0110","0110","0101","0000","0000","0001","0011","0011","0011","0011","0101","0110","0111","0111","0111","0100","0110","1000","0101","0011","0111","0101","0111","0111","0101","0011","0011","0010","0101","0110","0111","0111","0111","0110","0100","0011","0011","0110","0111","0111","0111","0111","0111","0101","0101","0101","0101","0100","0011","0011","0010","0001","0010","0011","0011","0011","0010","0010","0010","0001","0001","0010","0010","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0010","0001","0010","0011","0011","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0101","0101","0101","0100","0001","0001","0001","0001","0010","0011","0011","0010"),
("0101","0011","0011","0010","0010","0001","0001","0001","0011","0101","0110","0110","0100","0011","0011","0111","0111","0111","0100","0001","0001","0001","0001","0101","1000","0111","0110","0110","0111","0100","0000","0000","0000","0000","0010","0011","0010","0100","0101","0101","0101","0001","0000","0000","0000","0010","0100","0011","0010","0010","0001","0001","0110","0101","0011","0001","0000","0000","0000","0010","0100","0100","0011","0100","0100","0010","0001","0010","0001","0010","0010","0010","0001","0001","0000","0000","0000","0000","0010","0010","0011","0010","0100","0001","0000","0011","0001","0000","0010","0011","0001","0000","0000","0000","0000","0000","0001","0001","0000","0011","0100","0010","0001","0001","0001","0011","0011","0011","0011","0011","0011","0011","0011","0001","0000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0101","0011","0100","0100","0011","0101","0100","0011","0101","0011","0011","0101","0011","0100","0101","0011","0101","0100","0011","0100","0100","0100","0101","0101","0100","0110","0100","0101","0101","0100","0101","0100","0100","0100","0100","0100","0011","0010","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0100","0101","0110","0101","0110","0100","0010","0100","0011","0011","0011","0011","0011","0100","0100","0101","0101","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0011","0010","0001","0000","0000","0000","0010","0100","0000","0001","0001","0010","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0101","0101","0100","0100","0100","0101","0111","0101","0110","0100","0011","0001","0000","0000","0001","0011","0101","0110","0110","0110","0010","0000","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0010","0010","0010","0011","0100","0011","0100","0101","0101","0110","0110","0111","0111","0111","0101","0001","0000","0001","0011","0011","0011","0100","0110","0110","0111","0111","0110","0011","0101","0110","0011","0011","0110","0111","0111","0111","0101","0011","0011","0010","0110","0111","0111","0111","0111","0110","0100","0011","0011","0110","0111","0111","0111","0111","0111","0101","0101","0101","0101","0100","0011","0011","0010","0001","0001","0001","0010","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0001","0001","0010","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0001"),
("0001","0001","0001","0001","0001","0001","0001","0010","0010","0101","0110","0110","0100","0011","0011","0110","0111","0111","0101","0100","0100","0100","0100","0100","0111","0111","0111","0101","0110","0100","0010","0010","0010","0001","0100","0011","0001","0011","0100","0110","0110","0001","0001","0000","0000","0010","0100","0011","0100","0110","0101","0001","0010","0100","0100","0001","0000","0000","0000","0001","0101","0100","0010","0010","0010","0010","0010","0011","0001","0001","0010","0010","0010","0001","0000","0000","0001","0001","0010","0101","0001","0001","0100","0100","0001","0001","0001","0001","0010","0011","0001","0000","0001","0000","0000","0000","0000","0001","0000","0010","0010","0001","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0001","0001","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0011","0100","0011","0100","0100","0011","0100","0011","0011","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0011","0011","0100","0100","0011","0101","0011","0100","0101","0011","0101","0100","0011","0110","0011","0011","0010","0010","0011","0010","0100","0101","0011","0101","0100","0011","0101","0100","0011","0101","0011","0100","0101","0011","0101","0101","0011","0101","0101","0100","0101","0101","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0011","0100","0101","0101","0101","0101","0011","0001","0010","0010","0011","0011","0010","0010","0011","0010","0010","0011","0100","0100","0101","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0100","0011","0010","0001","0001","0001","0010","0011","0001","0010","0010","0011","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0101","0100","0100","0100","0011","0101","0111","0110","0101","0011","0010","0001","0000","0001","0011","0100","0100","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0110","0110","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0011","0100","0101","0110","0110","0011","0110","0110","0110","0110","0111","0111","0111","0111","0110","0001","0000","0010","0011","0011","0011","0100","0110","0110","0111","0111","0101","0010","0100","0110","0011","0100","0110","0111","0110","0110","0101","0011","0011","0011","0110","0111","0111","0111","0111","0111","0101","0011","0011","0110","0111","0111","0111","0111","0111","0101","0101","0101","0101","0100","0010","0001","0001","0001","0001","0001","0001","0011","0011","0011","0010","0010","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0010","0001","0001"),
("0000","0000","0001","0000","0000","0001","0001","0011","0010","0101","0110","0110","0100","0011","0010","0110","0111","0111","0111","0110","0101","0101","0101","0101","0101","0100","0101","0011","0110","0110","0100","0101","0100","0101","0110","0100","0001","0101","0110","0111","0110","0100","0100","0100","0010","0011","0101","0100","0100","0111","0110","0010","0000","0010","0010","0001","0000","0000","0001","0001","0010","0011","0010","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0000","0000","0001","0001","0001","0011","0010","0001","0101","0101","0010","0000","0011","0001","0001","0010","0001","0000","0001","0000","0001","0001","0001","0001","0000","0010","0001","0000","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0011","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0100","0010","0000","0001","0010","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0101","0100","0011","0101","0011","0100","0101","0011","0100","0101","0011","0101","0101","0011","0101","0101","0011","0110","0100","0100","0110","0100","0100","0110","0011","0101","0110","0100","0101","0101","0011","0100","0110","0110","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0101","0100","0100","0100","0100","0101","0100","0101","0111","0110","0101","0011","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0011","0010","0010","0101","0110","0110","0110","0110","0101","0101","0101","0101","0101","0100","0110","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0101","0110","0111","0111","0111","0100","0110","0111","0110","0111","0111","0111","0111","0111","0110","0000","0000","0010","0011","0011","0011","0100","0110","0110","0111","0111","0101","0010","0011","0110","0101","0101","0111","0110","0110","0110","0101","0100","0100","0011","0110","0111","0111","0111","0111","0111","0101","0011","0011","0110","0111","0111","0111","0111","0111","0101","0101","0101","0101","0011","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0011","0010","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0000","0000","0000","0000","0001","0100","0010","0001"),
("0000","0000","0001","0000","0000","0000","0001","0011","0011","0101","0110","0110","0100","0011","0010","0110","0111","0111","0111","0111","0111","0101","0100","0110","0110","0100","0101","0101","0101","0110","0101","0110","0101","0101","0101","0011","0001","0101","0111","1000","1000","0110","0101","0101","0101","0101","0100","0011","0100","0100","0101","0011","0001","0100","0011","0001","0001","0000","0000","0010","0011","0010","0010","0010","0100","0011","0010","0010","0001","0010","0010","0010","0011","0001","0000","0000","0000","0000","0010","0001","0011","0010","0100","0100","0010","0000","0001","0001","0001","0010","0001","0000","0000","0001","0010","0010","0001","0001","0000","0010","0010","0000","0000","0000","0100","0110","0110","0110","0110","0110","0110","0101","0101","0011","0001","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0101","0100","0100","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0000","0001","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0101","0011","0100","0101","0010","0100","0101","0011","0101","0100","0011","0100","0100","0101","0110","0100","0110","0110","0100","0110","0110","0101","0110","0101","0101","0110","0101","0100","0011","0101","0101","0101","0101","0101","0100","0101","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0010","0011","0011","0011","0010","0010","0010","0010","0011","0011","0100","0011","0101","0110","0101","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0001","0001","0101","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0011","0100","0100","0100","0100","0100","0011","0011","0100","0011","0011","0100","0101","0110","0111","0111","1000","1000","0111","0100","0110","0111","0110","0110","0111","0111","0111","0111","0110","0001","0000","0001","0011","0011","0011","0100","0110","0110","0111","0111","0101","0010","0100","0101","0101","0110","0110","0111","0111","0110","0101","0011","0100","0100","0110","0111","0111","0111","0111","0111","0101","0011","0011","0101","0111","0111","0111","0111","0111","0101","0101","0101","0101","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0010","0001","0001","0000","0001","0001","0010","0010","0001","0001","0001","0001","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0100","0100","0010"),
("0000","0000","0000","0000","0001","0001","0001","0010","0010","0101","0110","0110","0100","0011","0010","0110","0111","0111","0111","0111","0111","0110","0110","0101","0110","0111","0111","0111","0111","0110","0110","0110","0110","0101","0100","0010","0001","0101","0111","0111","0111","0110","0110","0110","0110","0101","0100","0100","0100","0101","0101","0101","0011","0010","0011","0001","0001","0000","0000","0001","0101","0001","0010","0010","0010","0010","0001","0010","0011","0011","0010","0010","0011","0010","0001","0001","0001","0001","0010","0000","0001","0010","0001","0010","0010","0000","0000","0001","0001","0010","0000","0001","0000","0000","0001","0001","0010","0011","0001","0010","0001","0000","0000","0001","0100","1000","1000","1001","1001","1001","1001","1000","1000","0100","0001","0110","1000","1000","1001","1001","1000","1000","1001","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0010","0000","0001","0011","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0100","0100","0011","0101","0100","0011","0101","0100","0011","0110","0100","0010","0011","0101","0100","0011","0110","0100","0011","0110","0100","0011","0110","0100","0011","0110","0101","0100","0110","0101","0100","0110","0110","0101","0110","0110","0101","0110","0110","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0001","0001","0001","0001","0010","0010","0100","0100","0101","0101","0100","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0101","0101","0101","0101","0110","0110","0101","0110","0101","0100","0110","0111","0111","0110","0010","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0110","0111","0111","0110","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0010","0100","0101","0101","0101","0101","0101","0100","0100","0101","0101","0101","0110","0110","0110","1000","1000","1000","1000","0100","0011","0101","0100","0010","0010","0011","0100","0100","0101","0100","0001","0000","0001","0011","0011","0011","0100","0110","0110","0111","0111","0110","0100","0101","0110","0110","0110","0110","0111","0111","0110","0110","0011","0011","0100","0110","0111","0111","0111","0111","0111","0101","0011","0011","0101","1000","0111","0111","0111","0111","0101","0101","0101","0011","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0000","0001","0001","0000","0001","0000","0001","0001","0010","0100","0100"),
("0000","0000","0000","0001","0001","0001","0000","0010","0011","0101","0110","0110","0100","0011","0010","0110","0111","0111","0110","0111","0111","0111","0111","0111","0101","0110","0111","0111","0110","0110","0101","0101","0101","0100","0011","0010","0010","0100","0111","0111","0111","0111","0110","0110","0110","0100","0100","0100","0101","0100","0100","0101","0110","0010","0001","0001","0000","0000","0000","0000","0010","0010","0010","0001","0011","0011","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0001","0011","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0010","0001","0000","0000","0000","0001","0001","0001","0010","0001","0100","0011","0000","0000","0000","0011","0101","0101","0110","0110","0110","0111","0111","0111","0011","0001","0101","0110","0110","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0000","0001","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0010","0100","0101","0101","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0101","0100","0100","0101","0101","0011","0101","0101","0011","0101","0101","0011","0101","0101","0011","0101","0101","0011","0100","0110","0011","0101","0110","0100","0101","0111","0100","0101","0110","0100","0101","0110","0101","0101","0110","0101","0101","0110","0101","0101","0101","0100","0101","0110","0110","0100","0011","0010","0100","0100","0101","0101","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0011","0001","0010","0011","0011","0010","0000","0011","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0110","0101","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0010","0010","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0010","0100","0110","0110","0101","0101","0101","0101","0101","0101","0101","0110","0111","0111","0111","1000","1000","0111","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0001","0000","0010","0011","0011","0011","0100","0110","0110","0111","0110","0110","0101","0101","0110","0110","0110","0110","0111","0111","0110","0101","0011","0011","0100","0110","0111","0111","0111","0111","0111","0100","0011","0011","0100","0111","0111","0111","0111","0111","0101","0101","0101","0010","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0000","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0000","0001","0001","0001","0001","0001","0001","0001","0010","0010","0100","0100"),
("0000","0000","0000","0000","0000","0001","0000","0010","0100","0100","0110","0110","0100","0011","0010","0110","0111","0110","0110","0110","0110","0111","0110","0111","0111","0100","0100","0111","0110","0101","0100","0110","0101","0011","0010","0010","0010","0101","0110","0101","0100","0101","0110","0101","0100","0010","0001","0001","0011","0010","0000","0010","0101","0011","0001","0001","0000","0001","0001","0001","0010","0010","0010","0010","0010","0011","0010","0010","0001","0010","0010","0001","0001","0010","0011","0011","0010","0001","0010","0100","0001","0010","0001","0001","0010","0001","0010","0010","0000","0010","0001","0001","0001","0001","0001","0000","0001","0001","0001","0101","0101","0010","0000","0000","0010","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0110","0110","0110","0101","0100","0101","0101","0101","0101","0101","0110","0110","0110","0111","0111","1000","1000","0111","0111","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","0111","0111","0111","0110","0100","0001","0010","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0010","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0100","0100","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0101","0011","0100","0101","0011","0100","0101","0011","0100","0101","0011","0100","0110","0011","0100","0110","0100","0011","0011","0011","0100","0011","0100","0101","0011","0101","0101","0011","0101","0101","0011","0101","0101","0011","0101","0101","0100","0101","0101","0100","0101","0101","0100","0101","0101","0100","0101","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0001","0001","0001","0001","0000","0001","0001","0001","0000","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0010","0011","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0011","0100","0111","0111","0110","0101","0010","0101","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","0111","0111","0111","0101","0011","0010","0001","0001","0010","0010","0010","0011","0011","0010","0011","0011","0101","0101","0001","0000","0001","0011","0011","0011","0100","0110","0110","0110","0111","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0101","0011","0011","0100","0110","0111","0111","0111","0111","0111","0100","0010","0011","0011","0100","0110","0111","0111","0111","0100","0100","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0000","0001","0010","0010","0010","0010"),
("0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0011","0101","0100","0011","0010","0101","0110","0110","0110","0110","0110","0101","0110","0110","0101","0110","0101","0101","0101","0101","0100","0011","0100","0100","0010","0011","0010","0101","0101","0100","0100","0101","0101","0011","0100","0010","0011","0100","0010","0010","0010","0001","0010","0010","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0011","0001","0001","0010","0010","0001","0010","0010","0101","0010","0001","0011","0000","0001","0001","0001","0011","0001","0001","0001","0001","0001","0001","0001","0000","0001","0000","0001","0101","0101","0001","0000","0001","0010","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0101","0100","0110","0111","0101","0110","0111","0111","0111","0110","0101","0110","0111","0100","0100","0110","0101","0100","0101","0100","0101","0101","0100","0101","0100","0100","0110","0110","0101","0101","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0110","0110","0110","0110","0110","0101","0110","0110","0110","0110","0110","0111","0111","0111","0111","1000","0111","0111","1001","1001","1001","1001","1001","1001","1001","1001","1001","0101","0001","0010","0110","0111","1000","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0101","0010","0101","0101","0101","0101","0100","0100","0100","0100","0011","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0101","0101","0101","0010","0001","0001","0001","0001","0010","0001","0001","0010","0001","0001","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0011","0001","0100","0101","0101","0010","0001","0001","0010","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0010","0010","0011","0011","0011","0100","0011","0100","0100","0100","0100","0100","0011","0100","0100","0011","0101","0100","0011","0101","0100","0011","0101","0100","0011","0101","0100","0011","0101","0100","0011","0101","0100","0011","0101","0100","0011","0101","0100","0011","0101","0100","0100","0101","0100","0100","0101","0100","0100","0101","0100","0100","0101","0100","0100","0101","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0100","0001","0010","0100","0100","0100","0011","0001","0100","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0101","0011","0001","0001","0001","0010","0010","0010","0010","0001","0010","0011","0100","0100","0101","0110","0110","0001","0000","0010","0011","0011","0011","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0110","0101","0011","0011","0100","0111","0111","0111","0111","0111","0111","0101","0010","0011","0011","0110","0111","0111","0111","0111","0100","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0010","0001","0001","0010","0010","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001"),
("0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0010","0011","0010","0010","0101","0110","0101","0011","0010","0010","0011","0011","0011","0011","0100","0110","0101","0011","0100","0100","0011","0010","0010","0010","0010","0001","0010","0100","0011","0011","0100","0011","0010","0011","0011","0011","0101","0101","0101","0011","0011","0011","0010","0001","0000","0000","0000","0000","0000","0001","0001","0010","0010","0010","0011","0011","0001","0001","0001","0010","0010","0001","0000","0000","0001","0000","0010","0010","0010","0011","0001","0011","0001","0001","0000","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0010","0011","0001","0001","0001","0010","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0101","0101","0110","0110","0110","0111","0111","0111","0111","0110","0110","0110","0101","0110","0111","0110","0100","0101","0110","0101","0111","0111","0111","0111","0101","0101","0111","0110","0101","0101","0110","0100","0101","0101","0101","0111","0110","0111","0110","0101","0101","0111","0101","0100","0101","0111","0100","0100","0100","0101","0101","0101","0101","0101","0100","0100","0110","0110","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0100","0001","0010","0101","0100","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0111","1000","1000","1000","0111","0111","0111","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","0011","0111","1001","1001","1001","1000","1000","1000","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0011","0100","0101","0101","0101","0101","0011","0011","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0001","0010","0010","0010","0010","0011","0001","0100","0110","0110","0011","0010","0001","0011","0001","0001","0011","0000","0011","0010","0001","0011","0010","0001","0100","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0001","0000","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0101","0100","0011","0101","0100","0011","0101","0011","0011","0101","0011","0011","0110","0100","0011","0110","0011","0011","0100","0100","0101","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0000","0000","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0010","0001","0001","0010","0010","0010","0010","0010","0011","0100","0011","0100","0100","0100","0101","0111","0111","0110","0001","0000","0001","0011","0011","0011","0011","0110","0110","0111","0111","0111","0110","0110","0110","0110","0110","0111","0111","0111","0111","0110","0011","0011","0100","0111","0111","0111","0111","0111","0111","0101","0011","0011","0100","0110","0111","0111","0111","0111","0100","0010","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0000"),
("0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0010","0010","0001","0100","0110","0110","0011","0000","0000","0000","0000","0010","0100","0100","0100","0100","0101","0011","0001","0000","0000","0000","0001","0011","0001","0011","0011","0010","0010","0010","0001","0001","0010","0010","0011","0110","0110","0101","0101","0101","0101","0100","0001","0000","0000","0000","0000","0001","0100","0100","0100","0101","0011","0010","0011","0010","0010","0001","0000","0010","0011","0011","0010","0001","0001","0001","0010","0010","0110","0010","0010","0001","0001","0010","0001","0001","0010","0010","0010","0010","0001","0001","0000","0001","0001","0001","0001","0011","0001","0000","0000","0001","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0101","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0101","0101","0111","1000","0111","0100","0101","0101","0111","0111","0111","0111","0111","0111","0110","0101","0101","0111","0111","0101","0100","0110","0110","0110","0111","0111","1000","0111","0110","0110","0110","0101","0111","0111","0101","0100","0110","0101","0110","1000","0111","1000","0110","0101","0110","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0100","0101","0011","0001","0010","0101","0101","0110","0101","0100","0110","0101","0101","0110","0101","0100","0110","0111","0101","0101","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0111","0111","0111","0111","0110","0101","0110","0110","0110","0110","0110","0111","0111","0111","0111","1000","1001","1000","1000","1000","0011","0111","1001","1001","1001","1001","1001","1001","1001","1001","1000","0111","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","0110","0111","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0011","0100","0101","0101","0100","0011","0010","0011","0010","0010","0011","0010","0011","0010","0010","0010","0010","0001","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0010","0000","0010","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0101","0100","0011","0101","0100","0011","0110","0100","0011","0010","0100","0100","0011","0101","0100","0011","0110","0100","0011","0110","0101","0011","0110","0101","0011","0110","0101","0100","0110","0101","0100","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0100","0100","0100","0011","0100","0100","0110","0111","1000","0111","0110","0001","0000","0001","0010","0011","0010","0100","0110","0110","0111","0111","0111","0110","0110","0110","0111","0111","0111","0111","0111","0110","0101","0011","0011","0011","0110","0111","0111","0111","0111","0111","0101","0011","0011","0011","0110","0111","0110","0110","0111","0011","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0100","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0100","0011","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000"),
("0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0010","0001","0001","0100","0110","0101","0011","0000","0000","0000","0000","0011","0110","0100","0011","0101","0101","0011","0000","0000","0000","0000","0001","0100","0010","0010","0011","0001","0001","0000","0000","0000","0000","0000","0011","0101","0101","0100","0111","0101","0101","0101","0011","0001","0010","0000","0000","0001","0100","0100","0101","0100","0011","0011","0011","0010","0010","0001","0010","0011","0100","0011","0010","0001","0001","0001","0001","0001","0101","0100","0001","0000","0001","0010","0001","0000","0001","0001","0001","0001","0001","0010","0010","0001","0001","0000","0000","0011","0010","0001","0001","0001","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0100","0101","0110","0111","0111","0110","0110","0110","0111","0111","0110","0110","0111","0111","0101","0100","0101","0110","0111","0111","0111","0111","0111","0111","0110","0100","0110","1000","1000","0101","0100","0101","0111","0111","0111","0111","0111","0111","0111","0110","0110","0111","0111","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0001","0011","0101","0101","0111","0110","0110","0111","0111","0111","0111","0110","0101","0111","0110","0110","0110","0111","0101","0101","0110","0101","0110","0111","0111","0111","0110","0101","0111","0111","0101","0101","0111","0110","0100","0101","0100","0101","0101","0101","0101","0101","0100","0101","0111","0110","0110","0110","0101","0010","0100","0100","0100","0100","0100","0101","0101","0101","0101","0110","0101","1000","1001","1001","1001","1010","1010","1010","1010","1010","1010","0111","1000","1001","1010","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0000","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0011","0011","0010","0010","0010","0001","0011","0100","0011","0011","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0011","0101","0100","0011","0101","0100","0011","0101","0101","0011","0100","0101","0011","0100","0110","0011","0100","0101","0011","0100","0110","0011","0100","0110","0100","0100","0110","0100","0100","0110","0100","0100","0110","0101","0100","0110","0101","0100","0101","0101","0101","0101","0101","0100","0100","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0101","0100","0010","0011","0100","0100","0101","0111","0111","1000","0111","0110","0001","0000","0001","0011","0011","0011","0011","0110","0110","0111","0111","0111","0110","0110","0110","0111","0111","0111","0111","0110","0110","0101","0010","0010","0010","0011","0100","0111","0111","0111","0111","0101","0011","0011","0100","0111","0101","0011","0011","0110","0011","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0010","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0101","0100","0010","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0001","0000","0001","0000","0000"),
("0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0010","0001","0001","0100","0100","0011","0010","0000","0000","0000","0000","0010","0100","0101","0101","0100","0011","0010","0000","0000","0000","0000","0001","0100","0010","0001","0001","0010","0010","0000","0000","0000","0000","0000","0101","0100","0011","0101","0110","0101","0011","0101","0011","0010","0000","0000","0000","0001","0010","0011","0010","0011","0101","0110","0101","0010","0010","0001","0010","0001","0001","0000","0000","0001","0001","0001","0001","0000","0011","0110","0011","0000","0001","0010","0001","0000","0000","0000","0001","0000","0001","0010","0001","0001","0001","0001","0001","0010","0001","0000","0001","0001","0011","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0110","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","1000","0111","0101","0101","0110","0111","0111","0111","0110","0111","0111","1000","0110","0110","0111","0111","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0001","0010","0110","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0101","0101","1000","1000","0111","0100","0110","0110","0110","0111","0111","0111","0111","0110","0110","0110","0110","0111","1000","0111","0100","0110","0110","0110","0111","1000","1000","1000","0110","0101","0111","0111","0101","0110","0111","0110","0010","0100","0101","0110","0111","0110","0111","0110","0101","0101","0110","0101","0100","0101","0101","0101","0101","0110","0110","0110","0110","0110","0101","0110","0110","0110","0100","0101","0101","0101","0101","0110","0110","0110","0111","0111","0111","1000","1000","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","0111","0111","0111","0110","0110","0011","0000","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0100","0100","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0011","0101","0100","0011","0001","0001","0001","0000","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0101","0011","0100","0101","0011","0011","0101","0100","0011","0110","0100","0011","0101","0100","0011","0101","0101","0010","0100","0100","0011","0100","0110","0100","0100","0110","0100","0100","0101","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0011","0100","0100","0101","0111","1000","1000","0111","0110","0001","0000","0001","0010","0011","0011","0100","0110","0110","0111","0110","0110","0110","0110","0110","0111","0111","0111","0110","0110","0110","0101","0011","0010","0011","0011","0110","0111","0111","0111","0111","0101","0011","0011","0100","0111","0110","0100","0101","0110","0101","0100","0011","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0010","0011","0010","0010","0001","0001","0001","0001","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0101","0100","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0000","0001"),
("0000","0001","0000","0000","0000","0000","0001","0001","0000","0000","0001","0011","0010","0001","0001","0011","0101","0110","0011","0000","0000","0000","0000","0010","0100","0011","0100","0011","0010","0010","0001","0000","0001","0000","0000","0011","0010","0001","0011","0011","0011","0000","0000","0000","0000","0000","0100","0100","0100","0100","0011","0001","0001","0010","0010","0001","0001","0000","0000","0001","0100","0011","0010","0010","0011","0100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0001","0001","0100","0101","0001","0001","0011","0010","0001","0001","0010","0001","0000","0001","0001","0001","0000","0001","0001","0001","0001","0000","0001","0011","0001","0011","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0101","0101","0110","0100","0010","0010","0010","0010","0010","0011","0011","0101","0111","0111","0111","0111","0101","0110","0101","0101","0101","0101","0101","0110","0110","0110","0111","0111","0111","0111","0110","0110","0111","0111","0111","0110","0110","0111","0110","0110","0110","0110","0111","0111","0111","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0001","0010","0110","0101","0101","0110","0111","0111","0110","0110","0111","0111","0111","0110","0110","1000","1000","0111","0100","0101","0110","0111","0111","0111","0111","0111","0111","1000","0101","0101","1000","1000","1000","0100","0110","0110","0111","0111","1000","1000","1000","0111","0111","0110","0101","0111","1001","1000","0100","0010","0101","0111","0111","1000","1000","1000","0110","0110","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0110","1000","0011","0010","0011","0010","0011","0011","0011","0011","0011","0010","0010","0101","0110","0101","0110","0111","0011","0010","0011","0011","0011","0100","0100","0100","0100","0100","0101","0101","0110","0111","1000","1000","0111","0110","0111","0111","0111","0111","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","0100","0000","0100","0111","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0011","0100","0010","0000","0000","0000","0001","0010","0011","0100","0100","0100","0100","0100","0011","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0101","0011","0011","0101","0011","0011","0101","0011","0011","0101","0010","0011","0101","0011","0011","0100","0100","0100","0101","0101","0101","0010","0100","0100","0100","0101","0111","1000","0111","0111","0110","0001","0000","0001","0010","0011","0011","0100","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0110","0111","0111","0110","0101","0010","0011","0011","0100","0110","0111","0111","0111","0110","0100","0010","0011","0011","0110","0101","0101","0110","0110","0110","0110","0111","0110","0110","0100","0010","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0001","0001","0001","0010","0001","0001","0001","0001","0010","0011","0011","0011","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000"),
("0000","0000","0000","0000","0001","0000","0000","0001","0000","0000","0001","0011","0011","0010","0010","0100","0101","0101","0011","0000","0001","0001","0000","0010","0011","0100","0011","0010","0010","0010","0001","0001","0001","0000","0000","0010","0001","0001","0011","0101","0100","0001","0000","0000","0000","0000","0010","0011","0011","0010","0001","0010","0100","0011","0011","0001","0000","0000","0000","0000","0010","0011","0100","0101","0110","0101","0101","0011","0001","0000","0000","0000","0000","0000","0000","0001","0001","0000","0010","0011","0001","0001","0011","0001","0001","0010","0010","0000","0001","0010","0001","0001","0000","0000","0001","0000","0001","0001","0000","0000","0000","0001","0101","0010","0010","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0101","0101","0101","0011","0001","0001","0001","0001","0001","0001","0001","0010","0110","0111","0111","0110","0101","0101","0010","0000","0001","0001","0000","0001","0001","0001","0101","0110","0111","0111","0110","0101","0101","0011","0010","0011","0011","0011","0100","0100","0101","0110","0111","0111","0111","0101","0110","0111","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","1000","0101","0100","0101","0101","0101","0101","0101","0101","0101","0011","0001","0010","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1000","1000","0111","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1000","1000","1000","0100","0110","0110","1000","1000","0111","0111","0111","1000","1000","0110","0110","1000","1001","1000","0101","0010","0101","1000","1000","0111","0111","0111","0111","1000","0110","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0110","0111","0110","0011","0100","0100","0100","0100","0110","0110","0110","0101","0100","0100","0110","0110","0101","0101","0111","0100","0010","0100","0011","0011","0100","0100","0100","0100","0011","0011","0100","1000","0110","0101","0110","0111","0010","0010","0010","0010","0010","0011","0010","0011","0011","0011","0011","0101","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0011","0000","0011","0110","0101","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","0111","0111","0111","0111","0110","0110","0011","0010","0101","0100","0001","0000","0000","0000","0001","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0101","0101","0101","0101","0100","0011","0100","0101","0111","0111","0111","1000","1000","0111","0110","0100","0100","0101","0100","0011","0011","0011","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110","0100","0011","0011","0011","0100","0110","0110","0101","0101","0100","0011","0001","0001","0010","0011","0101","0110","0110","0110","0111","0111","0110","0110","0100","0011","0011","0011","0010","0010","0010","0010","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0011","0010","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0000","0001","0001","0001","0000","0000","0000","0001","0000","0000","0000","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0000","0001","0001","0000","0001","0001","0001","0001","0000","0000","0000","0001"),
("0000","0000","0000","0000","0001","0001","0001","0000","0000","0001","0010","0010","0010","0010","0001","0101","0110","0101","0010","0000","0000","0000","0000","0010","0011","0010","0010","0011","0011","0010","0000","0000","0000","0000","0000","0001","0001","0010","0100","0010","0011","0001","0000","0000","0000","0001","0011","0001","0001","0100","0100","0010","0010","0100","0100","0001","0000","0000","0000","0001","0010","0100","0110","0110","0101","0101","0100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0010","0000","0001","0001","0000","0011","0011","0000","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0000","0000","0000","0010","0100","0010","0010","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0101","0101","0101","0100","0001","0001","0001","0001","0001","0001","0001","0010","0101","0111","0111","0111","0100","0101","0010","0001","0001","0001","0001","0010","0001","0001","0100","0110","0111","0111","0110","0101","0100","0001","0000","0000","0000","0000","0000","0000","0001","0101","0110","0111","0111","0101","0101","0011","0000","0001","0001","0001","0010","0010","0010","0101","0110","0111","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0010","0101","0101","0110","0101","0101","0101","0110","0110","0110","0110","0110","0111","0111","1000","1000","0111","0101","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","1000","1000","1000","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1000","1001","1000","0101","0010","0101","0111","0111","0111","0110","0111","0111","0111","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0111","1000","0101","0011","0100","0101","0110","0111","0111","0111","0111","0111","0110","0101","0100","0100","0111","1000","0101","0011","0100","0101","0101","0110","0110","0110","0110","0111","0101","0101","0100","0110","0101","0111","0110","0110","0010","0100","0100","0100","0100","0101","0101","0101","0101","0011","0011","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0010","0000","0100","0101","0100","0101","0100","0100","0101","0100","0100","0100","0100","0100","0100","0110","0101","0101","0110","0110","0100","0101","0100","0100","0101","0101","0101","0101","0101","0101","0110","0110","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1000","0110","1000","1001","0111","0001","0010","0110","0101","0001","0000","0000","0000","0011","0110","0110","0111","0111","0111","0110","0110","0100","0101","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0101","0101","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0010","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0101","0101","0100","0101","0110","0101","0111","1001","1010","1000","0111","1000","1000","1000","0110","0100","0101","0111","0101","0010","0010","0011","0110","0110","0111","0111","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0101","0011","0011","0100","0101","0111","0100","0001","0001","0001","0001","0001","0001","0010","0100","0101","0110","0110","0110","0101","0100","0011","0011","0100","0100","0011","0011","0010","0001","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0000","0000","0000","0000","0001","0001"),
("0000","0001","0000","0000","0001","0001","0001","0000","0000","0001","0001","0001","0001","0010","0001","0011","0100","0100","0010","0001","0000","0000","0000","0001","0010","0010","0010","0100","0011","0010","0000","0000","0000","0000","0000","0001","0001","0010","0011","0010","0100","0010","0000","0000","0000","0000","0011","0100","0011","0100","0100","0010","0011","0100","0011","0000","0001","0001","0001","0001","0001","0100","0101","0100","0010","0011","0011","0010","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0011","0011","0000","0000","0001","0000","0011","0011","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0000","0000","0000","0010","0100","0011","0001","0100","0100","0100","0101","0101","0101","0100","0100","0011","0001","0101","0110","0110","0100","0010","0001","0010","0001","0001","0010","0001","0010","0110","0111","0111","0111","0101","0101","0010","0001","0001","0001","0001","0011","0001","0001","0100","0110","0111","0111","0110","0101","0101","0001","0001","0000","0000","0001","0001","0001","0001","0100","0110","0111","0111","0101","0101","0011","0000","0000","0000","0000","0001","0001","0000","0010","0110","0111","0111","0101","0100","0101","0101","0101","0101","0101","0101","0101","0011","0001","0010","0101","0101","0110","0010","0000","0000","0000","0001","0001","0001","0001","0101","0110","1000","1000","0111","0101","0110","0011","0010","0011","0011","0011","0011","0011","0100","0110","0111","1000","1000","1000","0110","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","0101","0010","0101","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0111","1000","0110","0100","0101","0110","0111","0111","0110","0110","0110","0110","0111","0110","0101","0100","1000","1000","0110","0100","0101","0101","0110","0111","0111","0111","0111","0111","0111","0111","0101","0100","0101","1000","0111","0100","0011","0100","0101","0110","0110","0111","0111","0111","0110","0101","0101","0100","0110","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0101","0111","0110","0101","0111","0111","0111","0111","0110","0101","0110","0111","0101","0101","0110","0111","0101","0110","0101","0101","0110","0110","0110","0110","0101","0100","0101","0111","0101","0101","0101","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0101","0110","0110","0101","0101","0101","0100","0010","0101","0110","0100","0000","0001","0001","0001","0001","0000","0001","0001","0100","0101","1001","1001","1001","1001","1001","1001","0111","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","0111","0110","0111","0110","0101","0100","0100","0101","0110","0110","0110","0101","0101","0110","0101","0100","0101","0101","0101","0101","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0010","0010","0100","0100","0100","0100","0011","0100","0011","0100","0011","0100","0100","0100","0100","0100","0110","1000","1001","1001","0110","1000","1000","0111","0111","0111","1000","1000","1000","0110","0100","0101","0111","0101","0010","0010","0011","0101","0110","0111","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0110","0100","0010","0011","0100","0100","0111","0101","0001","0000","0000","0000","0000","0001","0101","0110","0110","0101","0100","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0010","0000","0000","0000","0010","0011","0011","0011","0100","0011","0100","0011","0100","0100","0100","1000","0110","0010","0001","0001","0010","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0101","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0001","0000","0001","0001","0001","0000","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0000","0000","0000","0000","0001","0000"),
("0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0000","0000","0010","0010","0010","0100","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0100","0010","0001","0001","0000","0000","0000","0001","0000","0010","0011","0110","0101","0001","0000","0000","0000","0000","0011","0100","0110","0110","0011","0011","0011","0100","0010","0001","0001","0001","0001","0001","0000","0001","0010","0011","0010","0010","0011","0010","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0011","0101","0011","0001","0001","0000","0010","0010","0001","0001","0001","0001","0000","0001","0000","0000","0000","0001","0011","0001","0000","0000","0011","0101","0010","0001","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0101","0110","0101","0100","0010","0001","0010","0001","0010","0010","0001","0010","0110","0111","0111","0111","0101","0101","0010","0001","0001","0001","0001","0011","0001","0001","0100","0110","0111","0111","0110","0101","0101","0001","0001","0000","0000","0010","0010","0001","0000","0100","0110","0111","0111","0101","0101","0011","0000","0000","0001","0001","0010","0001","0000","0010","0110","0111","0111","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0001","0010","0101","0101","0101","0010","0000","0000","0000","0001","0010","0000","0000","0011","0110","0111","1000","0111","0101","0101","0001","0000","0001","0001","0000","0001","0001","0000","0011","0110","1000","1000","0111","0101","0110","0010","0001","0001","0001","0001","0010","0010","0010","0101","0111","1000","1000","1000","0110","0010","0100","0100","0101","0101","0101","0101","0110","0110","0111","0111","0111","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0111","1001","0110","0101","0110","0111","0111","0111","0111","0110","0110","0111","0110","0110","0110","0110","1000","1000","0110","0100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0110","1000","0111","0101","0100","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0100","0111","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0101","0110","0110","0111","0111","0111","0111","1000","0110","0110","0110","0101","0111","1000","1000","0101","0101","0110","0110","0110","1000","1000","1000","1000","0110","0110","0111","0110","0101","0110","0110","0111","0100","0110","0101","0110","0111","0111","0111","0111","0101","0101","0110","0111","0101","0101","0110","0111","0100","0101","0100","0100","0010","0010","0010","0010","0001","0000","0000","0000","0000","0001","0010","0011","0100","0110","0110","0111","0111","0111","0111","0110","0111","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1001","1001","1001","0111","0100","0100","0101","0110","0111","1000","1001","1001","1001","1000","1000","0100","0110","0110","0101","0011","0010","0100","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0100","0010","0010","0100","0100","0011","0011","0100","0100","0011","0011","0011","0100","0100","0100","0110","1000","1010","1001","1001","0110","0101","0101","0110","0110","0111","1000","1000","1000","1000","0110","0100","0101","0111","0101","0011","0011","0101","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0110","0100","0011","0011","0011","0011","0011","0101","0101","0001","0000","0001","0000","0000","0001","0011","0100","0011","0011","0011","0011","0011","0010","0011","0100","0011","0100","0100","0100","0100","0010","0001","0001","0001","0010","0011","0100","0100","0011","0010","0011","0011","0011","0011","0101","1011","1001","0001","0000","0000","0000","0011","0011","0100","0100","0100","0011","0011","0100","0100","0100","0100","0101","0101","0100","0100","0011","0011","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0000","0001","0001","0000","0000","0001","0001","0000","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001"),
("0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0011","0011","0010","0010","0001","0001","0001","0010","0010","0001","0001","0010","0011","0010","0010","0010","0010","0001","0001","0001","0000","0010","0011","0101","0100","0010","0010","0010","0001","0001","0100","0100","0110","0110","0100","0011","0011","0010","0010","0010","0000","0000","0001","0001","0010","0001","0001","0100","0011","0001","0001","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","0101","0100","0001","0001","0000","0001","0010","0000","0001","0010","0001","0000","0000","0000","0001","0001","0000","0010","0001","0001","0001","0010","0011","0010","0001","0100","0100","0100","0100","0100","0100","0100","0100","0011","0000","0101","0110","0101","0100","0001","0001","0001","0001","0001","0010","0001","0010","0101","0111","0111","0111","0101","0101","0010","0001","0001","0001","0001","0011","0001","0001","0100","0110","0111","0111","0110","0101","0101","0010","0001","0000","0000","0010","0010","0000","0001","0100","0110","0111","0111","0101","0101","0011","0000","0000","0001","0001","0010","0001","0000","0010","0110","0111","0111","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0001","0010","0101","0101","0110","0010","0000","0000","0000","0001","0010","0000","0000","0011","0110","0111","1000","0111","0101","0110","0010","0001","0001","0001","0001","0010","0001","0001","0011","0110","1000","1000","0111","0101","0110","0010","0001","0001","0001","0000","0010","0001","0001","0011","0110","1000","1000","1000","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0011","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0111","1001","0110","0101","0110","0101","0101","0101","0101","0101","0101","0110","0110","0110","0111","0111","1000","1000","0110","0101","0111","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","0111","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0111","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0100","0101","0110","0111","0111","0111","0111","0111","1000","1000","0110","0101","0111","1000","1000","0101","0100","0101","0111","0111","1000","0111","0111","0111","0111","0111","0101","0100","0111","1000","1000","0100","0101","0110","0110","0110","0111","0111","1000","0111","0110","0110","0110","0101","0110","0111","0111","0101","0101","0110","0101","0101","0110","0001","0001","0001","0010","0001","0000","0000","0000","0000","0000","0010","0100","0101","0100","0100","0100","0100","0100","0101","0110","0110","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0110","0110","0110","0110","0101","0110","0101","0101","0101","0011","0010","0011","0100","0011","0100","0110","0110","1000","1000","1000","1000","0011","0011","0011","0010","0010","0010","0100","0111","1001","1001","1010","1010","1010","1010","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","0111","0011","0100","0111","0111","0111","0111","0111","0110","0110","0110","0101","0101","0111","1000","1001","1001","0111","0101","0100","0101","0101","0101","0110","0110","0111","0111","1000","1000","1000","0110","0100","0101","0111","0101","0010","0010","0100","0101","0110","0111","0111","0110","0111","0111","0111","0111","0111","0110","0101","0100","0100","0101","0101","0101","0101","0101","0110","0110","0001","0001","0000","0000","0000","0001","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0100","0011","0001","0000","0001","0001","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0001","0000","0001","0001","0011","0011","0100","0100","0100","0100","0101","0101","0101","0100","0011","0011","0100","0100","0011","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0001","0000","0001","0001","0000","0000","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001"),
("0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0001","0000","0001","0010","0011","0011","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0010","0100","0101","0100","0011","0011","0011","0010","0010","0100","0101","0110","0100","0010","0001","0011","0011","0100","0001","0000","0000","0000","0001","0011","0001","0000","0011","0110","0011","0001","0001","0001","0000","0000","0001","0000","0000","0000","0000","0000","0000","0010","0100","0011","0100","0011","0000","0000","0000","0001","0000","0001","0011","0001","0001","0000","0001","0001","0001","0000","0001","0001","0001","0001","0010","0011","0001","0001","0100","0100","0100","0100","0100","0100","0100","0101","0011","0000","0101","0110","0101","0100","0000","0000","0000","0000","0000","0000","0000","0001","0101","0111","0111","0111","0101","0101","0010","0000","0001","0001","0001","0001","0001","0000","0011","0110","0111","0111","0110","0101","0101","0001","0001","0001","0001","0010","0010","0001","0001","0100","0110","0111","0111","0110","0101","0011","0001","0000","0001","0001","0010","0001","0000","0001","0101","0111","0111","0101","0100","0101","0101","0101","0101","0101","0101","0101","0011","0001","0010","0101","0101","0110","0010","0000","0000","0000","0001","0011","0000","0001","0011","0110","0111","1000","0111","0101","0110","0010","0001","0001","0001","0001","0010","0001","0001","0011","0110","0111","1000","0111","0101","0110","0010","0001","0001","0001","0001","0010","0001","0001","0011","0110","0111","1000","0111","0101","0010","0001","0001","0001","0001","0000","0001","0001","0001","0001","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","1001","0110","0100","0110","0010","0000","0001","0001","0001","0000","0001","0001","0001","0100","0110","1000","1000","0110","0101","0110","0110","0011","0011","0011","0011","0011","0011","0100","0100","0101","0111","0111","1000","0111","0101","0101","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","0111","1000","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0111","1000","1000","0101","0101","0110","0111","0111","0111","0110","0110","0111","0111","0111","0110","0101","1000","1000","1000","0101","0101","0101","0111","0111","0111","0111","0111","0111","0111","0111","0100","0101","0111","1000","0111","0100","0100","0101","0110","0111","0111","0100","0000","0000","0001","0001","0000","0010","0011","0000","0000","0001","0100","0100","0101","0101","0101","0101","0100","0100","0111","0111","0100","0110","0110","0101","0101","0111","0110","0110","0111","0101","0101","0110","0111","0101","0101","0101","0111","0100","0101","0100","0100","0100","0011","0011","0010","0011","0011","0010","0100","0100","0100","0100","0100","0011","0010","0010","0010","0001","0001","0010","0010","0011","0101","0110","0110","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1001","1001","1001","1001","1000","1000","0011","0100","1001","1001","1010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0110","0101","0110","0101","0110","0100","0101","0110","0110","0111","0111","0111","0111","1000","0111","0100","0101","0111","0101","0010","0010","0101","0111","0111","0111","0111","0111","0111","0111","0111","0110","0101","0101","0110","0110","0110","0110","0111","0111","0110","0111","0110","0100","0001","0001","0001","0001","0001","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0100","0100","0100","0010","0001","0001","0001","0101","0110","0011","0011","0011","0011","0100","0100","0100","0100","0011","0000","0000","0001","0001","0000","0001","0011","0100","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0001","0001","0000","0000","0010","0010","0010","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0000","0000","0000","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0000","0001","0001","0000","0000","0000","0001","0001","0010","0011","0010","0011","0010","0001","0001"),
("0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0010","0010","0001","0001","0001","0001","0001","0010","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0000","0010","0101","0110","0100","0011","0101","0110","0011","0101","0100","0100","0100","0011","0001","0101","0110","0100","0101","0001","0000","0001","0000","0001","0011","0101","0011","0000","0011","0011","0010","0010","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0010","0011","0100","0101","0001","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0000","0100","0100","0000","0001","0100","0100","0100","0100","0100","0101","0100","0101","0011","0000","0101","0110","0101","0100","0000","0000","0001","0000","0001","0001","0001","0010","0101","0111","0111","0111","0101","0101","0010","0000","0001","0001","0000","0001","0000","0000","0011","0110","0111","0111","0110","0101","0101","0001","0000","0000","0000","0000","0001","0001","0001","0100","0110","0111","0111","0101","0101","0011","0000","0001","0001","0001","0001","0001","0001","0010","0101","0111","0111","0101","0100","0100","0100","0101","0101","0101","0101","0101","0011","0001","0001","0101","0101","0110","0010","0000","0000","0000","0001","0010","0001","0000","0011","0110","0111","0111","0111","0101","0110","0010","0001","0001","0001","0001","0011","0001","0001","0011","0110","0111","1000","0111","0101","0110","0010","0001","0001","0001","0001","0010","0001","0001","0011","0111","1000","1000","1000","0101","0010","0011","0010","0001","0000","0000","0010","0001","0000","0001","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0110","0101","0100","0111","1001","0110","0100","0101","0010","0001","0001","0001","0000","0001","0010","0001","0001","0011","0110","1000","1000","0110","0100","0110","0100","0000","0000","0001","0001","0000","0001","0001","0000","0001","0101","0111","1000","0111","0101","0101","0111","0011","0001","0001","0001","0001","0010","0010","0010","0010","0101","0111","1000","0110","0100","0100","0101","0101","0100","0101","0101","0101","0101","0101","0011","0000","0100","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","1000","1000","1000","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","1000","1000","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0100","0001","0010","0110","0110","0110","0110","0011","0101","0111","0100","0010","0010","0100","0000","0000","0001","0010","0010","0101","0101","0101","0101","0100","0101","0111","0111","0101","0110","0110","0110","0110","0111","0111","0111","0111","0110","0110","0110","0101","0110","0111","0111","0101","0101","0110","0110","0110","1000","0111","0110","0100","0010","0011","0100","0111","0100","0010","0100","0101","0100","0010","0011","0011","0100","0001","0011","0010","0001","0001","0011","0101","0110","0101","0101","0110","0110","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0110","0110","0010","0011","0110","0110","0111","0111","0111","0111","0111","0111","1000","1000","0111","0110","0101","0110","1000","0111","0101","0110","0101","0101","0110","0110","0111","0111","0111","0111","1000","0110","0100","0100","0101","0011","0010","0010","0100","0110","0110","0110","0110","0110","0110","0101","0101","0101","0111","1000","1000","0111","0110","0111","0110","0101","0011","0010","0010","0010","0001","0001","0000","0001","0001","0001","0010","0011","0011","0011","0011","0100","0011","0011","0011","0100","0011","0011","0011","0100","0100","0010","0001","0001","0001","0011","0111","0101","0011","0100","0011","0100","0011","0011","0011","0010","0000","0000","0001","0001","0001","0001","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0100","0011","0001","0001","0001","0001","0011","0100","0011","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0000","0000","0001","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0000","0000","0000","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001"),
("0000","0001","0000","0001","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0010","0001","0011","0001","0000","0000","0001","0001","0010","0011","0010","0001","0001","0001","0010","0011","0010","0001","0010","0001","0001","0011","0100","0101","0100","0101","0101","0101","0100","0101","0011","0100","0100","0001","0011","0100","0011","0101","0100","0010","0000","0001","0001","0001","0100","0101","0100","0001","0000","0010","0110","0101","0100","0010","0001","0001","0010","0001","0001","0000","0000","0001","0001","0001","0010","0100","0011","0001","0000","0010","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0010","0001","0000","0001","0100","0010","0000","0001","0100","0100","0100","0101","0101","0101","0100","0100","0011","0001","0101","0110","0101","0100","0001","0001","0010","0001","0010","0010","0001","0010","0101","0111","0111","0111","0101","0101","0010","0001","0001","0010","0001","0010","0000","0000","0011","0110","0111","0111","0110","0101","0101","0001","0000","0000","0000","0001","0001","0000","0000","0100","0110","0111","0111","0101","0101","0011","0000","0000","0000","0000","0000","0000","0000","0001","0101","0111","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0101","0101","0110","0010","0000","0001","0001","0001","0001","0001","0001","0011","0110","0111","0111","0111","0101","0101","0010","0001","0001","0001","0001","0010","0001","0001","0011","0110","0111","0111","0111","0101","0110","0010","0001","0001","0001","0001","0010","0001","0001","0011","0110","0111","0110","0101","0010","0001","0010","0010","0001","0001","0001","0001","0001","0000","0001","0110","0110","0101","0101","0101","0110","0110","0110","0101","0101","0110","0101","0100","0111","1000","0110","0101","0101","0010","0001","0001","0000","0000","0010","0010","0001","0001","0011","0110","1000","1000","0110","0101","0101","0101","0001","0001","0001","0001","0001","0010","0001","0001","0001","0101","0110","1000","0111","0101","0100","0110","0010","0001","0001","0001","0001","0001","0001","0001","0001","0011","0111","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0101","0101","0010","0010","0010","0010","0010","0011","0011","0011","0101","0110","0111","1000","1000","0110","0110","0111","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","1000","1000","0101","0110","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0111","0111","0110","0011","0010","0000","0100","0100","0011","0101","0100","0101","0101","0100","0010","0011","0011","0000","0000","0000","0010","0100","0101","0101","0101","0101","0100","0101","1000","1000","0101","0101","0101","0111","0111","0111","0111","0111","0111","0111","0111","0100","0101","1000","1000","1000","0101","0101","0101","0110","0111","1000","0111","0111","0101","0011","0010","0100","0100","0110","0101","0100","0100","0010","0010","0100","0101","0101","0100","0101","0101","0010","0010","0010","0010","0100","0110","0110","0111","0110","0101","0110","0101","0110","0111","0110","0110","0111","0101","0101","0101","0101","0110","0011","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0110","0110","0111","1000","0111","0101","0111","0101","0101","0110","0110","0111","0111","0111","0111","1000","0110","0011","0011","0011","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0110","0110","0101","0110","0100","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0010","0100","0110","0101","0011","0011","0011","0001","0000","0000","0001","0010","0101","0111","0110","0011","0010","0011","0011","0011","0011","0010","0000","0000","0000","0001","0001","0001","0011","0011","0011","0011","0100","0011","0011","0011","0011","0100","0100","0100","0100","0101","0100","0010","0001","0001","0001","0011","0011","0100","0100","0100","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0000","0000","0001","0001","0001","0000","0000","0001","0000","0001","0001","0000","0001","0001","0000","0001","0001","0001","0001","0001","0000","0001","0001","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000"),
("0001","0001","0001","0000","0000","0001","0000","0001","0001","0000","0001","0000","0000","0000","0000","0000","0001","0010","0011","0001","0000","0001","0010","0001","0001","0001","0001","0001","0010","0001","0001","0010","0010","0001","0001","0001","0000","0010","0011","0100","0101","0110","0110","0100","0011","0101","0110","0100","0010","0010","0101","0100","0100","0110","0100","0010","0000","0000","0000","0000","0010","0010","0011","0010","0001","0001","0101","0101","0100","0001","0010","0010","0010","0010","0010","0000","0000","0001","0001","0001","0010","0010","0011","0001","0000","0010","0010","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0011","0010","0000","0000","0011","0010","0000","0001","0100","0100","0100","0100","0101","0101","0101","0100","0011","0001","0101","0110","0101","0100","0001","0001","0010","0001","0010","0010","0001","0010","0101","0111","0111","0111","0101","0101","0010","0001","0001","0001","0001","0011","0000","0000","0011","0110","0111","0111","0110","0101","0101","0010","0001","0000","0000","0010","0010","0000","0000","0100","0110","0111","0111","0110","0101","0011","0001","0000","0000","0000","0010","0001","0000","0001","0101","0111","0111","0101","0100","0101","0101","0101","0101","0101","0101","0101","0011","0001","0001","0101","0101","0110","0010","0000","0000","0000","0000","0001","0001","0000","0011","0110","0111","0111","0111","0101","0101","0010","0000","0000","0000","0000","0000","0000","0000","0010","0110","0111","0111","0111","0101","0110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0100","0100","0100","0011","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0111","1000","0110","0101","0101","0011","0001","0001","0000","0000","0010","0010","0000","0001","0011","0110","0111","1000","0110","0101","0110","0101","0001","0001","0001","0001","0001","0010","0001","0000","0001","0101","0110","1000","0111","0101","0100","0110","0011","0001","0001","0001","0001","0001","0010","0001","0001","0010","0111","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0101","0101","0000","0000","0000","0000","0000","0000","0000","0000","0011","0101","0111","1000","1000","0101","0101","0100","0000","0000","0000","0001","0001","0001","0001","0001","0101","0110","0111","0111","0111","0101","0110","0101","0100","0100","0100","0101","0101","0101","0101","0110","0101","0101","0111","0111","0111","0011","0010","0000","0010","0110","0011","0000","0001","0001","0010","0110","0011","0000","0010","0010","0001","0000","0010","0011","0100","0101","0101","0101","0100","0101","1000","1000","0101","0101","0101","0110","0110","0110","0101","0101","0110","0111","0110","0110","0110","0111","1000","1000","0101","0101","0110","0111","1000","0111","0111","0101","0111","0110","0100","0011","0100","0111","1000","0110","0100","0010","0011","0101","0111","0110","0101","0110","0100","0101","0100","0010","0010","0101","1000","1000","0111","0100","0101","0101","0110","0110","0111","0111","0111","0111","0101","0110","0111","0110","0110","0011","0010","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0110","0110","0110","0111","1000","0111","0101","0111","0101","0101","0110","0110","0111","0111","0111","0111","0111","0111","0011","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0101","0100","0100","0100","0100","0101","0101","0101","0100","0101","0100","0101","0100","0100","0100","0011","0101","0110","0101","0100","0100","0010","0010","0010","0001","0010","0011","0101","0111","0110","0011","0011","0011","0011","0100","0011","0001","0001","0001","0001","0000","0001","0001","0011","0100","0011","0011","0011","0011","0100","0011","0100","0011","0100","0100","0100","0100","0010","0001","0001","0001","0011","0100","0011","0100","0100","0101","0100","0011","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000"),
("0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0001","0001","0010","0011","0011","0001","0001","0010","0001","0010","0001","0010","0010","0001","0001","0001","0000","0001","0001","0001","0001","0001","0000","0010","0011","0100","0101","0101","0101","0010","0101","0110","0101","0011","0100","0011","0101","0011","0101","0110","0100","0010","0000","0000","0000","0000","0010","0001","0010","0011","0010","0000","0001","0011","0010","0011","0011","0011","0011","0100","0011","0001","0000","0010","0010","0001","0001","0000","0001","0000","0001","0000","0001","0000","0000","0010","0001","0000","0000","0000","0000","0000","0000","0011","0010","0000","0000","0000","0000","0001","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0000","0101","0110","0101","0100","0001","0010","0010","0001","0010","0010","0001","0001","0101","0111","0111","0111","0101","0101","0011","0001","0001","0001","0001","0011","0000","0000","0011","0110","0111","0111","0110","0101","0101","0010","0001","0001","0001","0010","0010","0000","0000","0100","0110","0111","0111","0110","0101","0100","0001","0000","0000","0000","0011","0001","0000","0001","0101","0111","0111","0101","0100","0101","0101","0101","0101","0101","0101","0101","0011","0001","0001","0101","0101","0110","0010","0000","0000","0000","0001","0011","0001","0000","0011","0110","0111","0111","0111","0101","0101","0010","0001","0001","0001","0000","0001","0000","0000","0010","0110","1000","0111","0110","0100","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","1000","1000","0101","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0011","0100","0101","0100","0011","0101","0011","0001","0001","0001","0000","0010","0010","0000","0001","0011","0110","0111","1000","0110","0100","0110","0101","0001","0010","0001","0001","0001","0010","0001","0000","0001","0101","0110","0111","0111","0101","0100","0110","0011","0001","0001","0001","0001","0001","0010","0001","0001","0010","0111","1000","0111","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0110","0101","0001","0000","0000","0000","0001","0001","0000","0000","0010","0101","0111","0111","1000","0101","0101","0100","0000","0000","0000","0000","0001","0001","0000","0000","0011","0110","0111","0111","0111","0101","0101","0011","0000","0000","0000","0000","0001","0001","0000","0000","0100","0100","0110","0111","0111","0010","0000","0000","0001","0001","0001","0000","0001","0001","0001","0011","0010","0010","0010","0011","0010","0001","0001","0010","0011","0101","0101","0100","0100","0101","1000","1000","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0111","1000","1000","0101","0101","0101","0101","0110","0110","0101","0011","0101","0110","0110","0110","0110","1000","1000","1000","0100","0011","0100","0100","0110","0101","0100","0101","0100","0110","0110","0010","0010","0100","1000","1000","1000","0100","0101","0110","0111","0111","0111","0111","0111","0111","0111","0111","0101","0101","0111","0011","0010","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0110","0110","0110","0111","0110","0111","0110","0111","0100","0101","0110","0110","0111","0111","0111","0111","0111","0101","0010","0001","0001","0001","0001","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0011","0011","0100","0100","0100","0100","0100","0100","0011","0100","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0100","0101","0100","0100","0100","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0001","0001","0001","0001","0010","0011","0100","0100","0100","0100","0101","0101","0100","0011","0011","0001","0000","0000","0000","0001","0001","0001","0000","0001","0001","0000","0000","0000","0000","0000","0001","0001","0000","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000"),
("0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0010","0000","0001","0001","0011","0010","0010","0011","0001","0001","0010","0001","0001","0000","0001","0001","0000","0000","0000","0010","0010","0011","0110","0110","0011","0110","0110","0101","0011","0100","0010","0010","0011","0100","0101","0101","0100","0001","0000","0000","0001","0001","0010","0011","0100","0010","0000","0000","0000","0000","0001","0010","0010","0011","0011","0010","0011","0011","0000","0001","0010","0011","0010","0000","0000","0000","0000","0001","0001","0000","0001","0010","0001","0000","0010","0101","0100","0001","0001","0011","0001","0000","0001","0000","0000","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0000","0101","0110","0110","0100","0001","0001","0001","0001","0010","0010","0000","0001","0110","0111","0111","0111","0101","0101","0011","0001","0001","0001","0001","0011","0000","0000","0011","0110","0110","0111","0110","0101","0101","0010","0001","0001","0001","0010","0010","0000","0000","0100","0110","0111","0111","0101","0101","0100","0001","0000","0000","0000","0011","0001","0000","0001","0101","0111","0111","0101","0100","0101","0101","0101","0101","0101","0101","0101","0011","0001","0001","0101","0101","0110","0011","0001","0000","0001","0001","0100","0001","0000","0011","0110","0111","0111","0111","0101","0101","0010","0001","0001","0001","0001","0011","0000","0000","0010","0101","0101","0011","0010","0010","0010","0011","0011","0100","0100","0100","0100","0011","0100","0100","0011","0010","0011","0101","1000","0110","0010","0010","0100","0100","0100","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0011","0101","0010","0000","0000","0001","0000","0001","0001","0001","0000","0011","0110","0111","1000","0110","0101","0101","0101","0001","0001","0001","0001","0001","0010","0001","0000","0001","0101","0110","0111","0111","0101","0100","0110","0011","0001","0001","0001","0000","0001","0010","0001","0000","0010","0111","1000","0111","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0110","0101","0001","0000","0000","0000","0001","0001","0000","0000","0010","0110","0111","0111","0111","0101","0101","0100","0001","0000","0000","0000","0010","0001","0000","0000","0011","0110","0111","0111","0111","0101","0101","0011","0000","0000","0000","0000","0010","0001","0000","0000","0100","0101","0010","0100","0111","0100","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0100","0001","0000","0001","0001","0010","0101","0101","0101","0011","0100","0100","0100","1000","1000","0101","0110","0101","0100","0100","0100","0101","0101","0101","0101","0110","0110","0110","0111","1000","1000","0110","0110","0111","0110","0111","0111","0110","0111","0110","0111","0110","0110","0110","1000","0111","0110","0101","0100","0010","0001","0100","0100","0011","0011","0100","0101","0011","0010","0010","0100","0111","1000","1000","0101","0101","0110","0110","0110","0110","0101","0101","0110","0111","0110","0110","0110","0110","0011","0010","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0111","1000","0111","0110","0111","0101","0101","0110","0110","0111","0111","0111","0111","0111","0100","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0001","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0100","0100","0100","0011","0100","0100","0011","0100","0100","0011","0011","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0001","0001","0001","0000","0001","0000","0001","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0001","0001","0001","0001","0000","0001","0001","0001","0001","0000","0001","0000","0001","0000","0001","0001","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","0001","0001"),
("0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0000","0000","0001","0000","0000","0000","0001","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0000","0001","0010","0001","0000","0000","0001","0001","0011","0101","0011","0100","0111","0101","0100","0100","0100","0011","0110","0101","0101","0101","0111","0100","0001","0000","0000","0001","0001","0011","0110","0101","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0001","0000","0000","0001","0001","0000","0000","0001","0000","0001","0100","0110","0101","0010","0000","0001","0001","0000","0010","0010","0000","0001","0001","0100","0100","0100","0100","0100","0101","0101","0101","0011","0000","0100","0101","0011","0011","0010","0010","0010","0011","0011","0011","0010","0010","0100","0110","0110","0110","0101","0101","0011","0001","0000","0001","0001","0011","0000","0000","0011","0110","0110","0111","0110","0101","0101","0010","0001","0001","0001","0010","0010","0000","0000","0100","0110","0111","0111","0101","0101","0100","0001","0000","0000","0000","0011","0001","0000","0001","0101","0111","0111","0101","0100","0101","0101","0101","0101","0101","0101","0101","0011","0001","0001","0101","0101","0110","0011","0001","0000","0001","0001","0100","0001","0000","0011","0110","0111","0111","0111","0101","0101","0010","0001","0001","0000","0000","0011","0001","0001","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0100","0100","0011","0100","0100","0100","0011","0010","0010","0010","0011","0001","0010","0011","0100","0100","0100","0011","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0011","0011","0100","0011","0011","0011","0010","0010","0011","0101","0110","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0110","0111","0111","0110","0101","0101","0101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0110","0111","0111","0101","0100","0110","0011","0000","0001","0001","0001","0001","0010","0001","0001","0010","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0110","0101","0001","0000","0000","0000","0001","0001","0000","0000","0010","0110","0111","0111","0111","0101","0101","0100","0001","0000","0000","0000","0010","0001","0000","0000","0011","0110","0111","0111","0111","0101","0110","0011","0000","0000","0000","0000","0010","0001","0000","0000","0100","0110","0010","0000","0001","0011","0101","0010","0000","0000","0000","0000","0001","0000","0000","0000","0010","0011","0000","0000","0001","0001","0001","0101","0101","0100","0011","0100","0100","0100","0111","1000","0101","0101","0011","0000","0000","0000","0000","0001","0001","0000","0001","0100","0101","0111","1000","1000","0110","0110","0011","0010","0010","0010","0011","0011","0011","0011","0100","0110","0110","1000","1000","0111","0101","0110","0011","0001","0100","0011","0010","0100","0100","0011","0011","0010","0011","0100","0101","0111","0111","0110","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0011","0010","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","0110","0110","0110","0111","0110","0100","0101","0111","0100","0101","0110","0110","0111","0111","0111","0111","0110","0010","0010","0001","0001","0001","0010","0011","0011","0010","0010","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0101","0100","0100","0100","0101","0101","0100","0100","0011","0011","0100","0100","0011","0100","0011","0001","0000","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0010","0001","0000"),
("0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0010","0011","0011","0011","0101","0100","0100","0011","0100","0010","0100","0110","0100","0100","0100","0101","0101","0010","0000","0000","0000","0000","0100","0110","0110","0100","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0011","0011","0000","0000","0001","0100","0100","0100","0100","0101","0100","0100","0100","0011","0001","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0010","0010","0110","0101","0101","0010","0001","0001","0010","0001","0011","0001","0001","0011","0110","0110","0111","0110","0101","0101","0010","0010","0001","0001","0010","0011","0001","0001","0100","0110","0110","0111","0101","0101","0100","0001","0000","0000","0000","0011","0001","0000","0001","0101","0111","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0101","0101","0110","0011","0001","0000","0001","0001","0100","0001","0000","0011","0101","0111","0111","0111","0101","0101","0010","0000","0000","0001","0010","0011","0011","0100","0100","0011","0100","0100","0100","0100","0011","0100","0101","0100","0100","0011","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0100","0100","0100","0100","0011","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0011","0010","0010","0001","0001","0100","0111","0101","0101","0011","0001","0001","0000","0001","0010","0010","0001","0001","0011","0110","0111","0111","0110","0101","0101","0101","0001","0001","0001","0000","0000","0001","0000","0000","0000","0100","0110","0111","0111","0101","0100","0110","0011","0000","0000","0000","0000","0000","0000","0000","0000","0010","0111","0111","0110","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0011","0000","0100","0110","0101","0101","0001","0001","0001","0001","0001","0001","0001","0001","0010","0101","0110","0111","0111","0101","0101","0100","0001","0000","0000","0000","0011","0010","0000","0000","0011","0110","0111","0111","0111","0101","0101","0011","0000","0000","0000","0000","0010","0010","0000","0000","0100","0110","0110","0010","0000","0000","0011","0000","0000","0000","0000","0000","0001","0001","0000","0000","0010","0010","0000","0000","0010","0010","0000","0010","0010","0010","0011","0100","0100","0100","0110","0111","0101","0101","0011","0000","0000","0000","0000","0010","0001","0000","0000","0011","0101","0111","0111","1000","0101","0101","0011","0001","0001","0001","0000","0000","0000","0000","0000","0011","0101","0111","0111","1000","0110","0100","0010","0001","0001","0001","0001","0010","0010","0010","0001","0010","0010","0011","0100","0110","0100","0100","0110","0101","0100","0100","0101","0101","0101","0101","0110","0110","0111","0111","0110","0011","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","0101","0110","0110","0110","0101","0101","0111","0101","0101","0110","0110","0111","0111","0111","0111","0101","0010","0011","0010","0010","0011","0010","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0001","0010","0010","0010","0010","0011","0011","0010","0001","0010","0001","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0100","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0010","0010","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0000","0001","0001","0001","0000","0001","0001","0000","0000","0001","0001","0000","0001","0001","0001","0010","0011","0010","0000","0001","0001","0000","0001","0001","0001","0001","0000","0000","0000","0001","0001","0000","0000","0000","0001","0001","0001","0010","0001","0001"),
("0000","0000","0000","0000","0000","0001","0000","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0001","0001","0000","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0010","0101","0001","0011","0101","0101","0100","0010","0100","0010","0100","0100","0011","0100","0011","0100","0100","0010","0001","0001","0001","0000","0101","0101","0100","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0010","0001","0000","0000","0000","0000","0000","0010","0010","0000","0000","0001","0000","0000","0011","0010","0000","0000","0001","0100","0100","0100","0100","0100","0101","0100","0010","0001","0010","0010","0010","0010","0011","0011","0011","0010","0011","0010","0011","0010","0010","0001","0011","0110","0111","0101","0110","0011","0001","0000","0000","0001","0011","0001","0000","0011","0110","0110","0111","0110","0101","0101","0010","0001","0001","0001","0001","0010","0001","0001","0100","0110","0111","0111","0101","0101","0100","0001","0010","0010","0010","0011","0010","0001","0010","0101","0111","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0101","0101","0110","0011","0001","0000","0001","0001","0100","0001","0000","0011","0110","0111","0111","0111","0101","0101","0010","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0011","0100","0011","0011","0011","0011","0011","0100","0011","0011","0100","0100","0100","0011","0100","0100","0100","0011","0011","0011","0011","0010","0010","0010","0001","0001","0001","0001","0001","0101","0111","0101","0101","0011","0001","0001","0001","0001","0010","0010","0001","0001","0011","0110","0111","0111","0110","0101","0101","0101","0001","0010","0001","0001","0001","0011","0001","0000","0001","0101","0110","0111","0111","0101","0100","0110","0011","0000","0000","0001","0000","0001","0001","0000","0000","0010","0110","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0110","0101","0001","0000","0000","0000","0001","0001","0001","0000","0010","0101","0110","0111","0111","0101","0101","0100","0001","0001","0001","0001","0010","0010","0001","0000","0011","0110","0111","0111","0111","0101","0101","0011","0001","0000","0001","0001","0010","0010","0000","0000","0100","0111","0100","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0001","0000","0001","0000","0001","0011","0011","0011","0101","0110","0111","0101","0110","0011","0000","0000","0000","0000","0010","0001","0000","0000","0011","0101","0110","0111","0111","0101","0100","0100","0010","0010","0001","0001","0001","0010","0010","0001","0010","0110","0111","0101","0110","0111","0011","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0100","0101","0100","0100","0110","0010","0000","0000","0000","0000","0000","0000","0000","0000","0100","0110","0110","0011","0010","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0110","0110","0110","0110","0110","0101","0101","0111","0100","0101","0110","0110","0111","0111","0111","0110","0011","0001","0001","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0100","0011","0100","0011","0011","0011","0010","0011","0011","0011","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0000","0001","0001","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0001","0001","0100","0101","0011","0000","0000","0000","0001","0010","0001","0001","0001","0000","0000","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001"),
("0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0010","0001","0000","0001","0010","0001","0000","0000","0000","0000","0000","0001","0001","0000","0001","0001","0010","0010","0010","0010","0001","0000","0001","0001","0000","0001","0011","0100","0001","0011","0011","0011","0100","0010","0010","0010","0100","0011","0100","0101","0101","0010","0001","0001","0001","0010","0001","0000","0100","0100","0100","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0010","0010","0010","0001","0000","0000","0000","0000","0010","0010","0000","0000","0000","0000","0000","0001","0000","0001","0010","0001","0100","0100","0100","0100","0101","0101","0100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0101","0111","0111","0101","0110","0011","0001","0001","0001","0001","0011","0001","0000","0011","0101","0110","0111","0110","0101","0101","0010","0001","0000","0000","0001","0010","0000","0000","0011","0110","0111","0111","0110","0101","0100","0001","0001","0001","0001","0010","0010","0001","0001","0101","0111","0111","0101","0100","0100","0101","0101","0101","0101","0101","0101","0011","0001","0001","0101","0101","0110","0011","0001","0010","0010","0001","0011","0010","0010","0011","0101","0111","0111","0111","0101","0101","0010","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0011","0101","0101","0110","0011","0001","0001","0000","0000","0010","0010","0000","0001","0011","0110","0111","0111","0110","0101","0101","0101","0001","0010","0001","0000","0001","0100","0001","0001","0001","0101","0110","0111","0111","0101","0100","0110","0011","0001","0000","0001","0000","0010","0010","0000","0000","0010","0110","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0110","0101","0001","0000","0000","0000","0001","0001","0000","0000","0010","0101","0110","0111","0111","0101","0101","0100","0000","0000","0000","0000","0000","0000","0000","0000","0011","0101","0111","0111","0111","0101","0101","0011","0000","0001","0001","0001","0001","0010","0001","0000","0001","0101","0100","0000","0010","0011","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0001","0000","0000","0000","0000","0001","0010","0010","0001","0000","0100","0101","0110","0101","0110","0011","0001","0000","0000","0000","0011","0010","0000","0000","0011","0101","0110","0111","0111","0101","0011","0010","0010","0010","0010","0001","0010","0010","0010","0001","0011","0110","0111","0110","0100","0101","0010","0010","0001","0011","0010","0001","0010","0010","0001","0001","0001","0010","0011","0100","0011","0101","0101","0100","0010","0000","0000","0001","0001","0001","0001","0000","0000","0011","0101","0110","0011","0010","0101","0101","0101","0101","0101","0100","0101","0101","0100","0100","0110","0110","0110","0110","0110","0101","0101","0111","0101","0101","0110","0101","0110","0111","0111","0101","0001","0001","0001","0010","0011","0011","0010","0010","0011","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0100","0100","0100","0100","0100","0100","0011","0100","0011","0011","0011","0100","0011","0011","0011","0010","0011","0100","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0011","0010","0001","0000","0001","0000","0001","0001","0000","0001","0000","0000","0001","0000","0000","0000","0001","0000","0010","0010","0001","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0001","0001","0001","0001","0010","0000"),
("0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0011","0011","0010","0001","0001","0001","0010","0001","0000","0000","0000","0000","0000","0001","0001","0000","0011","0100","0100","0010","0011","0011","0011","0001","0010","0010","0000","0001","0010","0001","0001","0001","0001","0001","0001","0000","0001","0010","0010","0010","0011","0011","0100","0010","0000","0000","0000","0000","0001","0010","0100","0100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0010","0010","0000","0000","0001","0000","0000","0000","0000","0001","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0011","0110","0111","0101","0110","0011","0001","0000","0000","0001","0011","0001","0000","0010","0101","0111","0111","0110","0101","0101","0010","0001","0000","0000","0010","0010","0000","0000","0011","0110","0111","0111","0110","0101","0100","0001","0001","0001","0000","0010","0001","0000","0001","0101","0111","0111","0101","0100","0101","0100","0100","0101","0101","0101","0101","0011","0001","0001","0101","0101","0110","0011","0001","0000","0000","0001","0011","0001","0001","0010","0101","0111","0111","0111","0101","0101","0010","0001","0001","0001","0001","0010","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0010","0011","0011","0100","0011","0001","0001","0000","0000","0010","0010","0000","0000","0010","0110","0111","0111","0110","0101","0101","0101","0010","0010","0001","0000","0001","0011","0010","0001","0001","0100","0110","0111","0111","0110","0100","0110","0011","0001","0000","0001","0000","0010","0011","0000","0000","0010","0110","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0110","0101","0001","0001","0001","0000","0001","0011","0000","0000","0010","0101","0110","0111","0111","0101","0101","0100","0000","0000","0000","0000","0001","0001","0000","0000","0011","0110","0111","0111","0111","0101","0101","0011","0000","0000","0000","0000","0010","0011","0001","0000","0000","0001","0101","0100","0010","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0011","0000","0001","0001","0000","0000","0010","0010","0000","0000","0000","0000","0010","0100","0101","0110","0011","0001","0001","0001","0000","0011","0010","0000","0000","0011","0101","0110","0111","0111","0110","0101","0010","0010","0010","0010","0010","0011","0010","0010","0010","0011","0110","1000","0110","0010","0011","0010","0010","0001","0001","0010","0010","0010","0010","0010","0001","0001","0010","0010","0011","0100","1000","0110","0101","0010","0001","0001","0001","0001","0001","0001","0000","0000","0010","0110","0111","0011","0010","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0110","0110","0110","0110","0110","0101","0101","0111","0100","0101","0110","0110","0111","0111","0110","0100","0001","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0000","0000","0000","0000","0001","0000","0000","0000","0001","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0001","0010","0001","0000"),
("0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","0001","0000","0000","0000","0000","0000","0000","0000","0010","0100","0101","0011","0100","0101","0100","0011","0010","0010","0000","0001","0000","0000","0000","0000","0000","0000","0000","0001","0011","0100","0011","0010","0011","0011","0100","0011","0001","0000","0000","0000","0001","0010","0010","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0010","0001","0001","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0010","0010","0000","0000","0001","0000","0000","0000","0000","0000","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0100","0011","0001","0000","0000","0000","0011","0001","0000","0010","0110","0111","0111","0110","0101","0101","0010","0010","0001","0000","0010","0010","0000","0000","0011","0110","0111","0111","0110","0101","0100","0001","0000","0000","0000","0011","0001","0000","0001","0101","0111","0111","0101","0100","0100","0100","0100","0101","0101","0101","0101","0011","0001","0001","0101","0101","0110","0011","0001","0000","0000","0001","0011","0001","0000","0010","0101","0111","0111","0111","0101","0101","0010","0001","0000","0000","0000","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0000","0000","0010","0110","0111","0111","0111","0101","0101","0101","0010","0010","0001","0000","0001","0100","0010","0010","0001","0100","0110","0111","0111","0101","0100","0110","0011","0001","0000","0001","0000","0010","0011","0000","0001","0010","0110","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0101","0101","0001","0001","0001","0000","0001","0011","0000","0000","0010","0101","0110","0111","0111","0101","0101","0100","0001","0000","0000","0000","0010","0010","0000","0000","0011","0101","0111","0111","0111","0101","0101","0011","0000","0000","0000","0001","0010","0010","0000","0000","0001","0001","0010","0100","0011","0011","0001","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0011","0011","0000","0001","0011","0001","0000","0001","0100","0010","0000","0000","0000","0000","0011","0101","0110","0011","0001","0001","0001","0001","0010","0001","0000","0000","0011","0101","0110","0111","0111","0110","0100","0010","0001","0010","0010","0010","0011","0010","0010","0011","0010","0101","0111","0111","0011","0010","0001","0011","0001","0000","0001","0001","0001","0010","0010","0001","0001","0010","0001","0011","0011","0101","0101","0101","0010","0001","0001","0001","0001","0001","0001","0001","0000","0010","0100","0100","0010","0010","0101","0101","0101","0101","0101","0100","0100","0011","0010","0101","0110","0110","0110","0110","0110","0101","0101","0111","0101","0101","0110","0110","0111","0111","0110","0011","0001","0010","0001","0010","0010","0010","0001","0001","0001","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0001","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0011","0010","0010","0010","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0000","0000","0000","0000","0001","0000","0000","0000","0001","0001","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0000"),
("0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0001","0100","0100","0011","0010","0010","0010","0011","0011","0001","0000","0000","0000","0011","0100","0011","0011","0101","0011","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0001","0000","0000","0010","0010","0000","0000","0001","0000","0000","0000","0001","0011","0000","0010","0100","0100","0100","0101","0100","0100","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0001","0000","0000","0000","0011","0001","0000","0010","0101","0110","0111","0110","0100","0101","0010","0010","0001","0000","0010","0011","0000","0000","0011","0110","0111","0111","0110","0101","0100","0001","0000","0000","0000","0011","0010","0000","0001","0101","0111","0111","0101","0101","0100","0101","0101","0101","0101","0101","0101","0100","0001","0001","0101","0101","0110","0011","0001","0000","0000","0000","0011","0000","0000","0010","0101","0111","0111","0111","0101","0101","0010","0001","0000","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0001","0011","0110","0111","1000","0111","0101","0101","0101","0010","0010","0010","0001","0001","0100","0010","0010","0001","0100","0110","1000","0111","0110","0100","0110","0011","0001","0000","0001","0000","0010","0011","0000","0000","0010","0110","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0101","0101","0001","0001","0000","0000","0001","0011","0000","0000","0010","0101","0110","0111","0111","0101","0101","0100","0001","0000","0000","0000","0010","0010","0000","0000","0011","0110","0111","0111","0111","0101","0101","0100","0000","0000","0001","0001","0010","0010","0001","0000","0011","0100","0000","0001","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","0100","0001","0001","0011","0001","0011","0011","0101","0101","0011","0001","0001","0001","0101","0101","0101","0011","0001","0000","0000","0001","0010","0000","0001","0000","0011","0101","0110","0111","0111","0101","0101","0011","0001","0010","0001","0001","0010","0010","0010","0010","0001","0010","0100","0110","0100","0010","0010","0011","0001","0001","0010","0010","0010","0010","0001","0010","0001","0010","0011","0011","0100","0100","0011","0100","0010","0001","0010","0010","0000","0001","0001","0010","0010","0010","0011","0011","0010","0010","0101","0101","0101","0101","0101","0100","0011","0100","0011","0100","0110","0110","0110","0110","0110","0101","0101","0111","0101","0101","0110","0110","0111","0111","0101","0010","0001","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0001","0010","0010","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","0011","0011","0100","0100","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0010","0011","0011","0011","0010","0001","0000","0000","0000","0001","0000","0000","0001","0001","0001","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000"),
("0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0100","0100","0101","0110","0100","0000","0000","0000","0001","0010","0100","0100","0011","0010","0010","0000","0000","0000","0001","0010","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0000","0001","0000","0001","0001","0001","0001","0001","0010","0010","0001","0000","0001","0011","0011","0000","0011","0100","0101","0100","0011","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0010","0011","0011","0011","0011","0100","0100","0100","0011","0010","0001","0001","0000","0011","0001","0000","0100","0110","0111","0111","0110","0101","0110","0010","0010","0001","0000","0010","0011","0000","0000","0011","0110","0111","0111","0110","0101","0100","0001","0000","0000","0000","0010","0010","0000","0001","0101","0111","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0101","0101","0101","0011","0001","0000","0000","0001","0011","0001","0000","0010","0101","0111","0111","0111","0101","0101","0010","0001","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0001","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0101","0101","0101","0101","0101","0100","0100","0011","0011","0001","0010","0110","0111","1000","0111","0101","0101","0101","0001","0010","0010","0010","0010","0011","0011","0011","0010","0101","0110","1000","0111","0101","0100","0110","0100","0001","0010","0010","0001","0010","0011","0000","0001","0010","0111","0111","0110","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0101","0101","0001","0001","0000","0000","0001","0011","0000","0000","0010","0101","0110","0111","0111","0101","0101","0100","0001","0000","0001","0000","0010","0010","0000","0000","0011","0110","0111","0111","0111","0101","0101","0011","0000","0000","0000","0000","0010","0010","0001","0000","0100","0110","0100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0110","0110","0010","0010","0100","0001","0010","0101","0101","0110","0100","0001","0100","0110","0111","0101","0100","0010","0001","0001","0000","0001","0010","0001","0001","0000","0010","0101","0110","0111","0111","0101","0101","0011","0000","0001","0001","0001","0001","0001","0001","0010","0001","0010","0100","0110","0100","0010","0010","0010","0010","0001","0001","0010","0001","0010","0001","0010","0010","0010","0001","0001","0011","0111","0011","0100","0011","0001","0010","0010","0001","0001","0001","0001","0001","0010","0011","0101","0011","0010","0101","0101","0100","0101","0100","0010","0010","0011","0011","0011","0100","0101","0101","0110","0110","0101","0101","0111","0101","0101","0110","0110","0111","0110","0011","0001","0010","0010","0010","0001","0001","0010","0011","0011","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0001","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0010","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0100","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0010","0001","0000","0000","0001","0001","0001","0000","0000","0001","0001","0001","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0000","0000","0000","0000","0001","0000","0000","0001","0001","0001","0000","0001","0010","0000","0000"),
("0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0010","0010","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0010","0010","0010","0010","0100","0100","0011","0001","0010","0011","0100","0101","0101","0101","0100","0011","0010","0001","0000","0000","0001","0010","0011","0011","0011","0011","0010","0001","0000","0001","0001","0001","0001","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0000","0001","0011","0100","0011","0100","0100","0011","0001","0001","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0011","0011","0011","0011","0100","0100","0011","0010","0010","0001","0010","0010","0010","0101","0110","0111","0111","0110","0110","0110","0010","0001","0001","0000","0001","0010","0000","0001","0110","0110","0111","0111","0110","0110","0101","0001","0000","0000","0000","0010","0001","0000","0001","0101","0111","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0101","0101","0101","0010","0001","0000","0000","0001","0011","0001","0000","0010","0101","0111","0111","0111","0101","0110","0010","0001","0010","0001","0001","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0100","0010","0010","0110","0111","1000","0111","0101","0101","0101","0001","0010","0001","0000","0000","0010","0001","0001","0001","0100","0110","1000","0111","0110","0100","0110","0100","0001","0010","0010","0010","0010","0011","0010","0010","0011","0111","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0110","0101","0001","0001","0001","0000","0001","0011","0000","0000","0010","0101","0110","0111","0111","0101","0101","0100","0001","0000","0000","0000","0010","0010","0000","0000","0011","0110","0111","0111","0111","0110","0110","0100","0010","0010","0001","0000","0000","0001","0010","0011","0100","0101","0101","0100","0100","0001","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0001","0101","0011","0000","0001","0011","0011","0100","0101","0100","0011","0010","0001","0100","0111","0111","0101","0101","0011","0010","0001","0000","0000","0010","0010","0000","0000","0010","0101","0110","0111","0111","0110","0101","0100","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0100","0111","0100","0011","0010","0011","0001","0001","0000","0010","0010","0001","0001","0010","0010","0010","0001","0010","0100","0111","0100","0011","0010","0001","0010","0001","0001","0001","0010","0001","0001","0011","0110","0111","0011","0001","0101","0101","0100","0100","0100","0011","0010","0011","0100","0011","0110","0101","0110","0110","0110","0101","0101","0111","0101","0101","0110","0110","0110","0110","0001","0001","0010","0010","0010","0010","0010","0011","0011","0010","0001","0001","0000","0010","0001","0001","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0010","0011","0011","0010","0011","0100","0100","0100","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0001","0001","0000","0001","0001","0001","0000","0000","0001","0001","0001","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0100","0100","0011","0001","0001","0000","0000"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0010","0100","0011","0001","0001","0010","0010","0010","0011","0100","0101","0100","0100","0011","0011","0011","0010","0010","0011","0100","0010","0000","0000","0001","0010","0010","0001","0001","0001","0001","0011","0010","0010","0001","0001","0001","0001","0001","0000","0001","0010","0000","0000","0000","0000","0000","0000","0001","0011","0100","0100","0011","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0100","0011","0011","0011","0011","0100","0100","0011","0011","0011","0010","0101","0101","0101","0101","0101","0111","0111","0111","0101","0101","0101","0100","0100","0100","0100","0100","0011","0011","0100","0110","0111","1000","0110","0101","0100","0010","0001","0010","0001","0001","0001","0001","0011","0110","0111","0111","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0001","0001","0101","0110","0111","0100","0001","0000","0000","0000","0011","0001","0000","0011","0110","0111","1000","0111","0100","0011","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0100","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0011","0011","0111","1000","0111","0101","0101","0101","0001","0010","0001","0000","0000","0011","0001","0001","0001","0100","0110","0111","0111","0110","0100","0110","0100","0001","0000","0000","0000","0010","0010","0000","0000","0010","0110","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0101","0101","0001","0010","0010","0010","0010","0011","0011","0011","0011","0101","0110","0111","0111","0101","0101","0100","0001","0010","0010","0001","0011","0011","0001","0001","0011","0110","0111","0111","0111","0101","0100","0011","0011","0100","0100","0011","0000","0000","0010","0010","0011","0011","0011","0100","0011","0010","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0001","0010","0000","0000","0000","0000","0010","0010","0010","0010","0000","0001","0001","0011","0101","0111","0101","0110","0100","0011","0001","0000","0000","0011","0010","0000","0000","0010","0101","0111","0111","0111","0110","0110","0100","0001","0010","0010","0001","0010","0010","0010","0001","0001","0010","0011","0100","0010","0010","0011","0010","0001","0001","0001","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0010","0100","0010","0001","0001","0001","0001","0001","0010","0001","0001","0011","0101","0110","0011","0001","0100","0100","0101","0100","0100","0100","0010","0011","0011","0011","0101","0110","0110","0110","0110","0101","0101","0111","0101","0101","0110","0101","0110","0100","0001","0001","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0010","0011","0100","0100","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0011","0010","0010","0001","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0010","0010","0010","0010","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0100","0100","0100","0011","0010","0010","0010","0010"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0010","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0000","0000","0001","0001","0010","0100","0011","0011","0010","0001","0010","0010","0010","0001","0010","0010","0001","0011","0011","0010","0001","0001","0001","0001","0001","0000","0001","0010","0000","0000","0000","0000","0000","0000","0010","0100","0100","0011","0001","0010","0010","0011","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0100","0100","0011","0100","0100","0100","0100","0011","0011","0011","0010","0011","0110","0110","0101","0101","0111","0111","0111","0101","0101","0110","0110","0110","0110","0101","0101","0101","0101","0101","0110","0111","1000","0110","0100","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0110","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0001","0001","0101","0101","0101","0100","0010","0010","0010","0010","0010","0001","0001","0101","0110","0111","0110","0011","0010","0010","0011","0100","0101","0101","0101","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0111","0111","0101","0101","0110","0001","0010","0001","0000","0000","0011","0001","0001","0001","0100","0110","1000","0111","0110","0100","0110","0011","0001","0000","0000","0000","0010","0011","0000","0001","0010","0110","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0100","0110","0101","0101","0010","0001","0000","0000","0001","0011","0000","0000","0010","0101","0110","0111","0111","0101","0101","0100","0001","0001","0010","0010","0010","0011","0010","0010","0011","0110","0111","0111","0110","0010","0010","0011","0011","0100","0100","0011","0010","0011","0001","0000","0000","0001","0010","0010","0010","0011","0100","0001","0001","0001","0000","0000","0000","0000","0000","0000","0010","0010","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0010","0111","0110","0110","0100","0011","0001","0001","0000","0011","0011","0000","0000","0011","0101","0111","0111","0111","0101","0110","0100","0000","0001","0010","0010","0011","0010","0010","0001","0001","0010","0010","0010","0010","0100","0100","0010","0000","0001","0001","0010","0001","0010","0010","0001","0001","0010","0011","0011","0010","0010","0011","0101","0011","0001","0001","0001","0001","0001","0001","0001","0000","0010","0110","0110","0011","0010","0100","0011","0100","0100","0011","0011","0011","0011","0011","0100","0101","0110","0110","0110","0110","0101","0101","0111","0101","0101","0101","0110","0110","0011","0001","0001","0010","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0011","0010","0010","0010","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0011","0100","0100","0100","0011","0100","0100","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0100","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0001","0010","0010","0010","0010","0010","0001","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0001","0000","0000","0000","0000","0000","0001","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0001","0010","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0011","0100","0101","0011","0011","0011","0010","0010","0010","0010","0001","0001","0010","0001","0001","0010","0011","0010","0001","0001","0001","0001","0001","0000","0001","0010","0000","0000","0000","0001","0000","0000","0010","0100","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0001","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0101","0111","0101","0110","0111","0111","0111","0101","0110","0111","1000","0111","0110","0110","0110","0111","0110","0101","0110","0111","0111","0111","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0111","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0001","0001","0101","0101","0100","0101","0101","0101","0101","0101","0100","0101","0101","0101","0100","0100","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0100","0101","0100","0100","0100","0101","0101","0100","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0011","0110","0110","0101","0110","0010","0010","0001","0001","0001","0011","0010","0001","0001","0100","0110","1000","0111","0110","0100","0110","0100","0001","0000","0000","0000","0010","0011","0000","0000","0001","0110","0111","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0011","0110","0101","0101","0010","0001","0000","0000","0001","0010","0000","0000","0001","0101","0110","0111","0111","0110","0101","0101","0001","0000","0000","0000","0010","0010","0000","0000","0010","0110","0111","0111","0111","0100","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0010","0011","0010","0001","0001","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0110","0110","0110","0011","0001","0001","0001","0000","0011","0011","0001","0001","0011","0110","0111","1000","0111","0100","0100","0100","0001","0001","0001","0010","0011","0001","0001","0001","0001","0010","0010","0010","0010","0100","0100","0011","0000","0001","0010","0010","0011","0010","0010","0001","0001","0010","0011","0010","0010","0011","0011","0011","0011","0001","0001","0010","0010","0010","0001","0000","0000","0010","0101","0110","0010","0001","0100","0101","0101","0011","0011","0011","0010","0010","0011","0100","0100","0101","0110","0101","0110","0101","0101","0111","0101","0101","0110","0101","0101","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0011","0100","0100","0011","0010","0010","0011","0011","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0100","0100","0100","0011","0011","0100","0011","0011","0011","0011","0010","0010","0010","0011","0011","0100","0100","0100","0011","0011","0010","0010","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0001","0001","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0011","0011","0100","0011","0100","0011","0011","0011"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0010","0001","0010","0010","0001","0010","0010","0011","0011","0010","0010","0001","0001","0001","0010","0011","0001","0000","0000","0001","0001","0011","0001","0010","0010","0010","0010","0011","0001","0000","0010","0100","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0110","0110","0110","0111","0111","0111","0101","0110","0111","1000","0111","0110","0110","0111","1000","0111","0110","0110","0111","0111","0110","0101","0110","0111","1000","0110","0110","0110","0111","1000","0110","0110","0111","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0101","0101","0101","0110","0110","0110","0101","0101","0101","0110","0110","0101","0010","0010","0011","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0010","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0011","0101","0101","0110","0010","0010","0001","0001","0001","0011","0010","0001","0001","0100","0110","1000","0111","0110","0100","0101","0100","0001","0000","0000","0000","0010","0011","0000","0000","0001","0110","0111","0110","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0011","0110","0101","0101","0010","0001","0000","0000","0001","0011","0000","0000","0001","0101","0110","0111","0111","0110","0101","0100","0001","0000","0000","0000","0010","0010","0000","0000","0010","0110","0110","0111","0111","0110","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0001","0010","0010","0100","0101","0110","0100","0010","0010","0001","0001","0011","0010","0011","0010","0011","0110","0110","0110","0101","0011","0100","0011","0001","0001","0000","0001","0001","0010","0001","0000","0001","0100","0011","0100","0010","0100","0101","0100","0001","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0101","0101","0010","0011","0010","0001","0001","0001","0010","0001","0001","0001","0000","0010","0101","0100","0010","0001","0011","0011","0100","0011","0011","0010","0010","0010","0010","0011","0100","0110","0110","0110","0101","0100","0101","0111","0101","0101","0110","0110","0011","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0011","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0010","0110","1000","1000","0100","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0000","0000","0001","0001","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0011","0011","0011","0100","0100","0100","0100","0100"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0010","0010","0010","0010","0001","0010","0010","0011","0011","0011","0011","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0011","0011","0010","0010","0001","0010","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0011","0010","0010","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0101","0110","0101","0110","0111","0111","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0111","0111","0111","0110","0101","0110","0111","0111","0111","0110","0110","0111","1000","0110","0110","0111","0111","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0101","0101","0101","0110","1000","0111","0110","0110","0110","1000","0110","0010","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0100","0011","0100","0100","0100","0011","0011","0011","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0011","0100","0100","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0011","0010","0100","0111","0111","0010","0001","0001","0001","0001","0011","0010","0001","0001","0101","0110","1000","0111","0110","0100","0110","0100","0001","0000","0000","0000","0010","0011","0000","0000","0001","0110","0111","0111","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0000","0100","0110","0101","0101","0010","0001","0001","0000","0001","0011","0000","0000","0001","0101","0110","0111","0111","0110","0101","0101","0001","0001","0000","0000","0010","0010","0000","0000","0010","0110","0110","0111","0111","0110","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0011","0001","0000","0001","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0001","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0011","0101","0010","0011","0100","0011","0001","0010","0010","0010","0011","0010","0010","0010","0011","0110","0110","0100","0100","0100","0100","0011","0001","0001","0001","0001","0001","0010","0010","0001","0010","0100","0100","0011","0100","0101","0100","0100","0001","0001","0010","0010","0010","0010","0010","0001","0010","0011","0010","0011","0101","1000","0011","0100","0010","0000","0000","0000","0000","0001","0001","0001","0000","0011","0101","0100","0010","0001","0011","0011","0100","0011","0010","0010","0001","0010","0011","0011","0100","0101","0101","0110","0100","0101","0101","0111","0100","0101","0110","0101","0010","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0100","0011","0011","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0111","1000","0111","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0101","0110","0110","0011","0011","0011","0011","0011","0100","0100","0010","0001","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0011","0011","0010","0010","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0010","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0011","0011","0011","0100","0100","0011","0100"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0100","0100","0100","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0001","0010","0010","0010","0011","0011","0010","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0001","0001","0011","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0001","0011","0011","0100","0100","0101","0111","0110","0100","0101","0110","0110","0110","0110","0110","0110","0110","0101","0101","0110","0111","1000","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0100","0101","0101","0110","0111","0111","0110","0110","0111","0101","0010","0011","0011","0100","0100","0100","0100","0011","0011","0100","0100","0100","0011","0100","0011","0100","0100","0011","0011","0100","0100","0011","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0101","0101","0011","0010","0010","0010","0010","0010","0001","0001","0010","0110","0110","1000","0111","0110","0101","0110","0101","0001","0000","0000","0001","0001","0010","0000","0000","0011","0111","0111","0111","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0011","0000","0011","0110","0101","0110","0010","0001","0001","0000","0001","0011","0000","0000","0001","0101","0110","0111","0111","0110","0101","0100","0001","0001","0001","0000","0010","0011","0000","0000","0010","0110","0101","0111","0110","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0001","0001","0001","0001","0000","0000","0000","0001","0001","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0011","0010","0010","0001","0010","0001","0010","0010","0010","0001","0010","0010","0010","0010","0011","0100","0011","0100","0011","0011","0010","0001","0001","0001","0001","0010","0010","0010","0001","0001","0010","0100","0100","0101","0100","0010","0011","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0110","0100","0100","0011","0011","0010","0000","0001","0001","0000","0001","0001","0000","0000","0010","0100","0011","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0100","0101","0101","0101","0110","0101","0101","0100","0100","0101","0011","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0101","0100","0100","0011","0011","0100","0100","0100","0100","0011","0001","0010","0010","0010","0010","0011","0100","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","1000","1010","1000","0010","0011","0011","0011","0011","0010","0011","0011","0010","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0100","0010","0010","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0001","0001","0000","0001","0001","0000","0000","0001","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0011","0011","0100","0100","0011","0011","0011"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0100","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0011","0011","0010","0010","0001","0010","0011","0011","0011","0100","0100","0011","0001","0010","0010","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0101","0101","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0101","0100","0011","0100","0100","0100","0101","0101","0101","0110","0110","0111","1000","1001","0110","0100","0100","0100","0100","0100","0100","0101","0101","0100","0001","0001","0101","0111","0110","0111","0111","0111","0111","0111","0101","0010","0010","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0101","1000","0111","0110","0011","0100","0100","0011","0011","0011","0011","0011","0010","0010","0010","0011","0110","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0011","0110","0110","0111","0010","0001","0001","0001","0001","0011","0001","0000","0010","0110","0110","0111","0111","0110","0110","0101","0010","0001","0001","0000","0010","0011","0000","0001","0011","0111","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0001","0001","0001","0010","0010","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0001","0001","0001","0001","0010","0010","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0001","0001","0001","0010","0010","0001","0001","0001","0010","0100","0011","0010","0011","0100","0100","0001","0010","0001","0001","0001","0010","0001","0010","0010","0001","0010","0100","0011","0010","0010","0011","0010","0001","0010","0001","0001","0010","0001","0001","0001","0010","0100","0011","0010","0010","0011","0011","0100","0011","0010","0011","0010","0010","0011","0010","0010","0100","0111","0101","0100","0101","0101","0100","0011","0011","0100","0011","0010","0001","0001","0001","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0010","0011","0101","0100","0011","0100","0100","0011","0010","0010","0010","0010","0011","0011","0010","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0011","0011","0010","0001","0011","0101","0110","0011","0010","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0011","0010","0011","1000","1001","0111","0010","0011","0011","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0011","0010","0010","0011","0011","0001","0001","0001","0010","0001","0001","0001","0001","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0011","0011","0100","0100","0011","0011","0011"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0100","0011","0011","0010","0010","0011","0011","0100","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0011","0010","0001","0001","0010","0011","0011","0011","0011","0100","0100","0011","0001","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0101","0101","0101","0100","0101","0101","0101","0101","0011","0001","0001","0001","0001","0001","0010","0001","0010","0001","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0101","0101","0101","0100","0100","0100","0011","0011","0011","0011","0011","0010","0010","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0001","0001","0011","0100","0011","0011","0100","0100","0101","0100","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0110","0110","0110","0101","0110","0110","0101","0110","0110","0110","0101","0110","1000","0111","0110","0011","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0110","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0011","0000","0011","0110","0100","0101","0011","0010","0010","0010","0010","0010","0010","0001","0011","0101","0110","0111","0111","0110","0110","0110","0010","0001","0001","0001","0010","0010","0000","0001","0100","0100","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0001","0001","0010","0010","0011","0010","0011","0001","0001","0000","0000","0001","0000","0000","0010","0010","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0001","0001","0010","0010","0001","0001","0001","0010","0001","0010","0010","0011","0010","0001","0010","0010","0010","0010","0001","0001","0001","0010","0010","0001","0010","0011","0110","0110","0011","0011","0011","0011","0001","0010","0010","0010","0010","0010","0001","0000","0001","0010","0010","0010","0011","0010","0010","0010","0010","0010","0001","0000","0001","0001","0001","0000","0001","0010","0011","0011","0010","0011","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0010","0100","0101","0100","0100","0100","0100","0100","0011","0011","0011","0010","0010","0010","0010","0010","0001","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0101","0101","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0011","0011","0001","0011","0011","0010","0001","0010","0011","0011","0010","0010","0010","0001","0001","0010","0010","0011","0011","0100","0100","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0010","0011","0011","0010","0101","1000","1000","0100","0010","0011","0011","0011","0100","0011","0011","0011","0011","0100","0011","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0001","0001","0000","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0000","0000","0000","0000","0001","0011","0011","0100","0100","0100","0100","0011","0011"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0011","0100","0100","0100","0101","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0001","0001","0010","0011","0011","0011","0011","0011","0100","0011","0011","0001","0010","0011","0100","0011","0100","0011","0011","0100","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0011","0001","0001","0010","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0101","0101","0101","0101","0100","0100","0100","0011","0011","0011","0101","0101","0101","0101","0101","0100","0011","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0011","0110","0111","1000","0111","0101","0101","0110","0111","1000","0111","0110","0110","1000","1000","0110","0100","0101","0110","0111","0111","0110","0101","0101","0110","0110","0110","0101","0110","1000","0111","0101","0101","0101","0101","0101","0100","0101","0101","0101","0101","0011","0000","0011","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0110","0111","0111","0110","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0010","0001","0000","0010","0100","0100","0100","0100","0011","0000","0000","0000","0000","0000","0000","0000","0010","0010","0001","0010","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0010","0010","0010","0010","0001","0001","0010","0010","0000","0001","0001","0001","0001","0010","0001","0001","0001","0010","0010","0001","0010","0110","0111","0101","0011","0011","0011","0010","0001","0010","0010","0010","0010","0001","0001","0001","0010","0001","0001","0011","0100","0010","0010","0001","0010","0010","0001","0000","0001","0010","0001","0000","0001","0010","0011","0001","0010","0010","0011","0011","0010","0010","0010","0010","0001","0010","0100","0011","0100","0011","0010","0010","0011","0011","0011","0100","0011","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0011","0011","0011","0100","0100","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0011","0011","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0010","0011","0011","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0010","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0100","0100","0011","0010","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0100","0100","0100","0100","0100","0011","0011"),
("0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0100","0100","0100","0011","0011","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0100","0100","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0100","0100","0101","0101","0101","0101","0011","0001","0001","0010","0100","0101","0101","0101","0100","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0100","0010","0100","0101","0110","0110","0110","0110","0100","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0101","0110","0111","0111","0101","0100","0101","0111","0111","0111","0110","0110","1000","1000","0111","0100","0101","0110","0111","1000","0111","0100","0101","0110","1000","0111","0110","0111","1000","0111","0101","0101","0101","0101","0101","0101","0100","0101","0100","0100","0011","0000","0100","0110","0101","0101","0110","0111","0110","0110","0110","0110","0110","0110","0110","0101","0110","1000","1000","0110","0101","0101","0110","0101","0110","0110","0110","0110","0101","0010","0010","0011","0010","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0010","0001","0001","0011","0011","0011","0010","0010","0000","0000","0000","0000","0000","0010","0001","0001","0000","0001","0001","0001","0001","0000","0000","0000","0000","0001","0010","0010","0001","0010","0011","0010","0001","0001","0000","0001","0010","0010","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0010","0101","0110","0011","0100","0011","0011","0010","0010","0010","0001","0001","0010","0010","0001","0001","0010","0011","0010","0011","0100","0010","0001","0010","0010","0010","0001","0001","0001","0010","0010","0001","0010","0010","0011","0010","0010","0010","0011","0010","0001","0010","0010","0001","0001","0011","0100","0011","0011","0011","0011","0011","0100","0010","0001","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0010","0011","0011","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0011","0100","0011","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0011","0011","0100","0011","0010","0011","0100","0011","0011","0011","0001","0010","0011","0011","0011","0011","0011","0011","0011","0011","0100","0011","0011","0100","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0100","0011","0011","0011","0010","0010","0001","0010","0011","0011","0011","0011","0100","0011","0011","0011","0011","0011","0011","0010","0010","0100","0100","0011","0010","0011","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0011","0100","0100","0100","0100","0100","0100","0011"),
("0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0010","0010","0001","0001","0010","0010","0010","0001","0010","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0010","0010","0010","0011","0011","0011","0011","0011","0011","0100","0100","0100","0010","0001","0011","0100","0100","0100","0100","0100","0100","0101","0101","0101","0100","0100","0101","0101","0101","0101","0011","0010","0001","0010","0011","0100","0101","0101","0100","0100","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0011","0100","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0010","0010","0010","0010","0011","0011","0011","0011","0010","0010","0010","0011","0010","0010","0011","0010","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0110","0110","0111","0110","0110","0110","0111","0110","0111","0110","0111","1000","1000","0111","0101","0101","0110","0111","0110","0111","0101","0101","0110","0111","0111","0110","0110","0111","0110","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0000","0011","0110","0101","0110","0110","1000","0111","0110","0110","0110","1000","1000","0110","0110","0111","0111","1000","0111","0101","0110","0111","0111","0110","0110","0110","0101","0010","0010","0011","0100","0001","0010","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0001","0001","0001","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0001","0001","0000","0001","0001","0001","0000","0001","0001","0000","0000","0000","0000","0010","0001","0001","0001","0011","0011","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0010","0001","0001","0001","0010","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0101","0101","0100","0101","0011","0010","0010","0010","0001","0001","0010","0001","0001","0001","0001","0010","0011","0001","0010","0010","0001","0001","0010","0010","0001","0001","0010","0010","0010","0010","0001","0001","0001","0010","0010","0010","0010","0010","0001","0010","0010","0010","0010","0011","0011","0100","0100","0100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0010","0010","0010","0011","0011","0010","0010","0011","0011","0011","0010","0011","0010","0010","0010","0010","0100","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0011","0011","0010","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0100","0011","0010","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100"),
("0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0010","0011","0011","0011","0011","0100","0011","0100","0100","0100","0100","0010","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0100","0100","0011","0010","0001","0010","0011","0100","0100","0101","0100","0100","0101","0101","0100","0100","0101","0101","0100","0100","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0100","0100","0101","0101","0100","0101","0101","0101","0100","0100","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0101","0100","0101","0101","0100","0100","0100","0011","0011","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0011","0011","0011","0010","0011","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0010","0011","0011","0100","0100","0100","0100","0100","0100","0100","0101","0110","0111","1000","1000","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0011","0000","0011","0101","0101","0110","0111","0111","0111","0110","0110","0110","0111","0111","0110","0110","0110","0111","0111","0110","0101","0110","0111","1001","0111","0110","0110","0010","0010","0011","0011","0011","0010","0000","0001","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0001","0001","0001","0001","0010","0010","0001","0001","0011","0010","0010","0010","0010","0011","0010","0010","0001","0001","0010","0010","0001","0001","0010","0001","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0011","0011","0011","0101","0011","0010","0001","0001","0010","0001","0001","0001","0001","0001","0010","0010","0011","0010","0010","0001","0001","0010","0010","0010","0001","0001","0010","0010","0010","0010","0001","0010","0001","0010","0010","0010","0010","0001","0001","0010","0010","0010","0010","0010","0010","0011","0100","0011","0010","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0001","0010","0010","0010","0010","0001","0010","0010","0010","0010","0010","0010","0011","0011","0011","0010","0010","0010","0010","0010","0011","0011","0100","0011","0011","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0101","0011","0100","0100","0011","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0100","0100","0100","0011","0011","0011","0011","0011","0011","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0001","0001","0001","0001","0000","0001","0001","0001","0010","0010","0001","0001","0000","0001","0001","0010","0010","0010","0011","0010","0010","0011","0011","0010","0010","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0100","0100")
);
begin
exctract:process (enable)
   begin
        if enable = '1' then
            data <= ROM(to_integer(unsigned(v_pos)), to_integer(unsigned(h_pos)));
            else data <= x"0";
        end if;
    end process;
end Behavioral;
